
module converter_out_I_n_node_interface_dut_ ( \n.buffer_full_in , 
        \n.receiving_data , \n.data_in , \n.buffer_full_out , \n.sending_data , 
        \n.data_out , buffer_full_out, sending_data, data_out, buffer_full_in, 
        receiving_data, data_in );
  input [15:0] \n.data_in ;
  output [15:0] \n.data_out ;
  output [15:0] data_out;
  input [15:0] data_in;
  input \n.buffer_full_in , \n.receiving_data , buffer_full_in, receiving_data;
  output \n.buffer_full_out , \n.sending_data , buffer_full_out, sending_data;


endmodule


module DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 ( 
        clk, rst_n, push_req_n, pop_req_n, diag_n, data_in, empty, 
        almost_empty, half_full, almost_full, full, error, data_out, peek_out
 );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] peek_out;
  input clk, rst_n, push_req_n, pop_req_n, diag_n;
  output empty, almost_empty, half_full, almost_full, full, error;


endmodule


module DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 ( 
        clk, rst_n, push_req_n, pop_req_n, diag_n, data_in, empty, 
        almost_empty, half_full, almost_full, full, error, data_out, peek_out
 );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] peek_out;
  input clk, rst_n, push_req_n, pop_req_n, diag_n;
  output empty, almost_empty, half_full, almost_full, full, error;


endmodule


module fifo_kev_63 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_127 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_63 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_127 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_126 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_63 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_126 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_63_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_63 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_63 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_63 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_63_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_62 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_125 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_62 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_125 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_124 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_62 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_124 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_62_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_62 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_62 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_62 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_62_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_61 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_123 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_61 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_123 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_122 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_61 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_122 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_61_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_61 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_61 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_61 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_61_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module converter_in_I_n_node_interface_dut__23 ( \n.buffer_full_in , 
        \n.receiving_data , \n.data_in , \n.buffer_full_out , \n.sending_data , 
        \n.data_out , buffer_full_out, sending_data, data_out, buffer_full_in, 
        receiving_data, data_in );
  input [15:0] \n.data_in ;
  output [15:0] \n.data_out ;
  output [15:0] data_out;
  input [15:0] data_in;
  input \n.buffer_full_in , \n.receiving_data , buffer_full_in, receiving_data;
  output \n.buffer_full_out , \n.sending_data , buffer_full_out, sending_data;
  wire   \n.buffer_full_in , \n.receiving_data , buffer_full_in,
         receiving_data;
  assign buffer_full_out = \n.buffer_full_in ;
  assign sending_data = \n.receiving_data ;
  assign data_out[15] = \n.data_in  [15];
  assign data_out[14] = \n.data_in  [14];
  assign data_out[13] = \n.data_in  [13];
  assign data_out[12] = \n.data_in  [12];
  assign data_out[11] = \n.data_in  [11];
  assign data_out[10] = \n.data_in  [10];
  assign data_out[9] = \n.data_in  [9];
  assign data_out[8] = \n.data_in  [8];
  assign data_out[7] = \n.data_in  [7];
  assign data_out[6] = \n.data_in  [6];
  assign data_out[5] = \n.data_in  [5];
  assign data_out[4] = \n.data_in  [4];
  assign data_out[3] = \n.data_in  [3];
  assign data_out[2] = \n.data_in  [2];
  assign data_out[1] = \n.data_in  [1];
  assign data_out[0] = \n.data_in  [0];
  assign \n.buffer_full_out  = buffer_full_in;
  assign \n.sending_data  = receiving_data;
  assign \n.data_out  [15] = data_in[15];
  assign \n.data_out  [14] = data_in[14];
  assign \n.data_out  [13] = data_in[13];
  assign \n.data_out  [12] = data_in[12];
  assign \n.data_out  [11] = data_in[11];
  assign \n.data_out  [10] = data_in[10];
  assign \n.data_out  [9] = data_in[9];
  assign \n.data_out  [8] = data_in[8];
  assign \n.data_out  [7] = data_in[7];
  assign \n.data_out  [6] = data_in[6];
  assign \n.data_out  [5] = data_in[5];
  assign \n.data_out  [4] = data_in[4];
  assign \n.data_out  [3] = data_in[3];
  assign \n.data_out  [2] = data_in[2];
  assign \n.data_out  [1] = data_in[1];
  assign \n.data_out  [0] = data_in[0];

endmodule


module flipflop_BITS2_23 ( clk, data_i, data_o );
  input [1:0] data_i;
  output [1:0] data_o;
  input clk;


  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS2_23 ( clk, enable_i, reset, data_i, data_o );
  input [1:0] data_i;
  input [1:0] data_o;
  input clk, enable_i, reset;
  wire   n10, n11, n1, n5, n7, n8, n9;
  wire   [1:0] write_data;

  AOI22X1 U5 ( .IN1(enable_i), .IN2(data_i[1]), .IN3(n10), .IN4(n1), .QN(n9)
         );
  AOI22X1 U6 ( .IN1(data_i[0]), .IN2(enable_i), .IN3(n11), .IN4(n1), .QN(n8)
         );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n9), .QN(write_data[1]) );
  NOR2X0 U4 ( .IN1(reset), .IN2(n8), .QN(write_data[0]) );
  AND2X1 U7 ( .IN1(data_o[1]), .IN2(n7), .Q(n10) );
  AND2X1 U8 ( .IN1(data_o[0]), .IN2(n5), .Q(n11) );
  flipflop_BITS2_23 FF ( .clk(clk), .data_i(write_data), .data_o({n7, n5}) );
endmodule


module flipflop_BITS1_87 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_87 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_87 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter2_23 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [1:0] request;
  output [1:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   tail_en, n1, n2;
  wire   [1:0] req_i;
  wire   [1:0] req_o;

  AND3X1 U10 ( .IN1(request[1]), .IN2(n1), .IN3(n2), .Q(grant[1]) );
  AND3X1 U11 ( .IN1(request[0]), .IN2(n2), .IN3(request[1]), .Q(tail_en) );
  INVX0 U6 ( .INP(request[0]), .ZN(n1) );
  NOR2X0 U7 ( .IN1(buffer_full_i), .IN2(n1), .QN(grant[0]) );
  INVX0 U8 ( .INP(buffer_full_i), .ZN(n2) );
  OA21X1 U9 ( .IN1(request[1]), .IN2(request[0]), .IN3(n2), .Q(grant_v_o) );
  register_BITS2_23 req_record ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i({1'b1, 1'b0}), .data_o({1'b0, 1'b0}) );
  register_BITS1_87 tail ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i(1'b1), .data_o(1'b0) );
endmodule


module flipflop_BITS2_22 ( clk, data_i, data_o );
  input [1:0] data_i;
  output [1:0] data_o;
  input clk;


  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS2_22 ( clk, enable_i, reset, data_i, data_o );
  input [1:0] data_i;
  input [1:0] data_o;
  input clk, enable_i, reset;
  wire   n10, n11, n1, n5, n7, n8, n9;
  wire   [1:0] write_data;

  AOI22X1 U5 ( .IN1(enable_i), .IN2(data_i[1]), .IN3(n10), .IN4(n1), .QN(n9)
         );
  AOI22X1 U6 ( .IN1(data_i[0]), .IN2(enable_i), .IN3(n11), .IN4(n1), .QN(n8)
         );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n9), .QN(write_data[1]) );
  NOR2X0 U4 ( .IN1(reset), .IN2(n8), .QN(write_data[0]) );
  AND2X1 U7 ( .IN1(data_o[1]), .IN2(n7), .Q(n10) );
  AND2X1 U8 ( .IN1(data_o[0]), .IN2(n5), .Q(n11) );
  flipflop_BITS2_22 FF ( .clk(clk), .data_i(write_data), .data_o({n7, n5}) );
endmodule


module flipflop_BITS1_86 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_86 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_86 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter2_22 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [1:0] request;
  output [1:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   tail_en, n1, n2;
  wire   [1:0] req_i;
  wire   [1:0] req_o;

  AND3X1 U10 ( .IN1(request[1]), .IN2(n1), .IN3(n2), .Q(grant[1]) );
  AND3X1 U11 ( .IN1(request[0]), .IN2(n2), .IN3(request[1]), .Q(tail_en) );
  INVX0 U6 ( .INP(request[0]), .ZN(n1) );
  NOR2X0 U7 ( .IN1(buffer_full_i), .IN2(n1), .QN(grant[0]) );
  INVX0 U8 ( .INP(buffer_full_i), .ZN(n2) );
  OA21X1 U9 ( .IN1(request[1]), .IN2(request[0]), .IN3(n2), .Q(grant_v_o) );
  register_BITS2_22 req_record ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i({1'b1, 1'b0}), .data_o({1'b0, 1'b0}) );
  register_BITS1_86 tail ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i(1'b1), .data_o(1'b0) );
endmodule


module dccl_63 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_62 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_61 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module controller3_nw ( clk, rst, .packet_addr({\packet_addr[2][7] , 
        \packet_addr[2][6] , \packet_addr[2][5] , \packet_addr[2][4] , 
        \packet_addr[2][3] , \packet_addr[2][2] , \packet_addr[2][1] , 
        \packet_addr[2][0] , \packet_addr[1][7] , \packet_addr[1][6] , 
        \packet_addr[1][5] , \packet_addr[1][4] , \packet_addr[1][3] , 
        \packet_addr[1][2] , \packet_addr[1][1] , \packet_addr[1][0] , 
        \packet_addr[0][7] , \packet_addr[0][6] , \packet_addr[0][5] , 
        \packet_addr[0][4] , \packet_addr[0][3] , \packet_addr[0][2] , 
        \packet_addr[0][1] , \packet_addr[0][0] }), local_addr, packet_valid, 
        buffer_full_in, grant_1, grant_2, grant_v, pop_v );
  input [7:0] local_addr;
  input [2:0] packet_valid;
  input [2:0] buffer_full_in;
  output [1:0] grant_1;
  output [1:0] grant_2;
  output [2:0] grant_v;
  output [2:0] pop_v;
  input clk, rst, \packet_addr[2][7] , \packet_addr[2][6] ,
         \packet_addr[2][5] , \packet_addr[2][4] , \packet_addr[2][3] ,
         \packet_addr[2][2] , \packet_addr[2][1] , \packet_addr[2][0] ,
         \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] ,
         \packet_addr[1][4] , \packet_addr[1][3] , \packet_addr[1][2] ,
         \packet_addr[1][1] , \packet_addr[1][0] , \packet_addr[0][7] ,
         \packet_addr[0][6] , \packet_addr[0][5] , \packet_addr[0][4] ,
         \packet_addr[0][3] , \packet_addr[0][2] , \packet_addr[0][1] ,
         \packet_addr[0][0] ;
  wire   \grant_2[1] , \request[2][1] , \request[2][0] , \request[1][1] ,
         \request[1][0] , \request[0][0] , n1;
  assign pop_v[1] = \grant_2[1] ;
  assign grant_2[1] = \grant_2[1] ;

  OR2X1 U3 ( .IN1(grant_v[0]), .IN2(grant_1[1]), .Q(pop_v[2]) );
  OR2X1 U4 ( .IN1(grant_1[0]), .IN2(grant_2[0]), .Q(pop_v[0]) );
  NOR2X0 U1 ( .IN1(n1), .IN2(buffer_full_in[0]), .QN(grant_v[0]) );
  INVX0 U2 ( .INP(\request[0][0] ), .ZN(n1) );
  arbiter2_23 arbiter_e ( .clk(clk), .rst(rst), .request({\request[1][1] , 
        \request[1][0] }), .buffer_full_i(buffer_full_in[1]), .grant(grant_1), 
        .grant_v_o(grant_v[1]) );
  arbiter2_22 arbiter_l ( .clk(clk), .rst(rst), .request({\request[2][1] , 
        \request[2][0] }), .buffer_full_i(buffer_full_in[2]), .grant({
        \grant_2[1] , grant_2[0]}), .grant_v_o(grant_v[2]) );
  dccl_63 dccl_s ( .packet_addr_y_i({\packet_addr[0][3] , \packet_addr[0][2] , 
        \packet_addr[0][1] , \packet_addr[0][0] }), .packet_addr_x_i({
        \packet_addr[0][7] , \packet_addr[0][6] , \packet_addr[0][5] , 
        \packet_addr[0][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[0]), 
        .east_req(\request[1][0] ), .local_req(\request[2][0] ) );
  dccl_62 dccl_e ( .packet_addr_y_i({\packet_addr[1][3] , \packet_addr[1][2] , 
        \packet_addr[1][1] , \packet_addr[1][0] }), .packet_addr_x_i({
        \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] , 
        \packet_addr[1][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[1]), 
        .local_req(\request[2][1] ) );
  dccl_61 dccl_l ( .packet_addr_y_i({\packet_addr[2][3] , \packet_addr[2][2] , 
        \packet_addr[2][1] , \packet_addr[2][0] }), .packet_addr_x_i({
        \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] , 
        \packet_addr[2][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[2]), 
        .east_req(\request[1][1] ), .south_req(\request[0][0] ) );
endmodule


module mux2_1_23 ( data0, data1, select0, select1, data_o );
  input [15:0] data0;
  input [15:0] data1;
  output [15:0] data_o;
  input select0, select1;
  wire   n1, n4, n5;

  AO22X1 U4 ( .IN1(data1[9]), .IN2(n5), .IN3(data0[9]), .IN4(n4), .Q(data_o[9]) );
  AO22X1 U5 ( .IN1(data1[8]), .IN2(n5), .IN3(data0[8]), .IN4(n4), .Q(data_o[8]) );
  AO22X1 U6 ( .IN1(data1[7]), .IN2(n5), .IN3(data0[7]), .IN4(n4), .Q(data_o[7]) );
  AO22X1 U7 ( .IN1(data1[6]), .IN2(n5), .IN3(data0[6]), .IN4(n4), .Q(data_o[6]) );
  AO22X1 U8 ( .IN1(data1[5]), .IN2(n5), .IN3(data0[5]), .IN4(n4), .Q(data_o[5]) );
  AO22X1 U9 ( .IN1(data1[4]), .IN2(n5), .IN3(data0[4]), .IN4(n4), .Q(data_o[4]) );
  AO22X1 U10 ( .IN1(data1[3]), .IN2(n5), .IN3(data0[3]), .IN4(n4), .Q(
        data_o[3]) );
  AO22X1 U11 ( .IN1(data1[2]), .IN2(n5), .IN3(data0[2]), .IN4(n4), .Q(
        data_o[2]) );
  AO22X1 U12 ( .IN1(data1[1]), .IN2(n5), .IN3(data0[1]), .IN4(n4), .Q(
        data_o[1]) );
  AO22X1 U13 ( .IN1(data1[15]), .IN2(n5), .IN3(data0[15]), .IN4(n4), .Q(
        data_o[15]) );
  AO22X1 U14 ( .IN1(data1[14]), .IN2(n5), .IN3(data0[14]), .IN4(n4), .Q(
        data_o[14]) );
  AO22X1 U15 ( .IN1(data1[13]), .IN2(n5), .IN3(data0[13]), .IN4(n4), .Q(
        data_o[13]) );
  AO22X1 U16 ( .IN1(data1[12]), .IN2(n5), .IN3(data0[12]), .IN4(n4), .Q(
        data_o[12]) );
  AO22X1 U17 ( .IN1(data1[11]), .IN2(n5), .IN3(data0[11]), .IN4(n4), .Q(
        data_o[11]) );
  AO22X1 U18 ( .IN1(data1[10]), .IN2(n5), .IN3(data0[10]), .IN4(n4), .Q(
        data_o[10]) );
  AO22X1 U19 ( .IN1(data1[0]), .IN2(n5), .IN3(data0[0]), .IN4(n4), .Q(
        data_o[0]) );
  INVX0 U2 ( .INP(select1), .ZN(n1) );
  AND2X1 U3 ( .IN1(select0), .IN2(n1), .Q(n4) );
  NOR2X0 U20 ( .IN1(n1), .IN2(select0), .QN(n5) );
endmodule


module mux2_1_22 ( data0, data1, select0, select1, data_o );
  input [15:0] data0;
  input [15:0] data1;
  output [15:0] data_o;
  input select0, select1;
  wire   n1, n4, n5;

  AO22X1 U4 ( .IN1(data1[9]), .IN2(n5), .IN3(data0[9]), .IN4(n4), .Q(data_o[9]) );
  AO22X1 U5 ( .IN1(data1[8]), .IN2(n5), .IN3(data0[8]), .IN4(n4), .Q(data_o[8]) );
  AO22X1 U6 ( .IN1(data1[7]), .IN2(n5), .IN3(data0[7]), .IN4(n4), .Q(data_o[7]) );
  AO22X1 U7 ( .IN1(data1[6]), .IN2(n5), .IN3(data0[6]), .IN4(n4), .Q(data_o[6]) );
  AO22X1 U8 ( .IN1(data1[5]), .IN2(n5), .IN3(data0[5]), .IN4(n4), .Q(data_o[5]) );
  AO22X1 U9 ( .IN1(data1[4]), .IN2(n5), .IN3(data0[4]), .IN4(n4), .Q(data_o[4]) );
  AO22X1 U10 ( .IN1(data1[3]), .IN2(n5), .IN3(data0[3]), .IN4(n4), .Q(
        data_o[3]) );
  AO22X1 U11 ( .IN1(data1[2]), .IN2(n5), .IN3(data0[2]), .IN4(n4), .Q(
        data_o[2]) );
  AO22X1 U12 ( .IN1(data1[1]), .IN2(n5), .IN3(data0[1]), .IN4(n4), .Q(
        data_o[1]) );
  AO22X1 U13 ( .IN1(data1[15]), .IN2(n5), .IN3(data0[15]), .IN4(n4), .Q(
        data_o[15]) );
  AO22X1 U14 ( .IN1(data1[14]), .IN2(n5), .IN3(data0[14]), .IN4(n4), .Q(
        data_o[14]) );
  AO22X1 U15 ( .IN1(data1[13]), .IN2(n5), .IN3(data0[13]), .IN4(n4), .Q(
        data_o[13]) );
  AO22X1 U16 ( .IN1(data1[12]), .IN2(n5), .IN3(data0[12]), .IN4(n4), .Q(
        data_o[12]) );
  AO22X1 U17 ( .IN1(data1[11]), .IN2(n5), .IN3(data0[11]), .IN4(n4), .Q(
        data_o[11]) );
  AO22X1 U18 ( .IN1(data1[10]), .IN2(n5), .IN3(data0[10]), .IN4(n4), .Q(
        data_o[10]) );
  AO22X1 U19 ( .IN1(data1[0]), .IN2(n5), .IN3(data0[0]), .IN4(n4), .Q(
        data_o[0]) );
  INVX0 U2 ( .INP(select1), .ZN(n1) );
  AND2X1 U3 ( .IN1(select0), .IN2(n1), .Q(n4) );
  NOR2X0 U20 ( .IN1(n1), .IN2(select0), .QN(n5) );
endmodule



    module node3_NODE_X0_NODE_Y0I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__ ( 
        \clk.clk , \reset.reset , \local_node.clk , 
        \local_node.buffer_full_in , \local_node.buffer_full_out , 
        \local_node.receiving_data , \local_node.sending_data , 
        \local_node.data_in , \local_node.data_out , \node_0.clk , 
        \node_0.buffer_full_in , \node_0.buffer_full_out , 
        \node_0.receiving_data , \node_0.sending_data , \node_0.data_in , 
        \node_0.data_out , \node_1.clk , \node_1.buffer_full_in , 
        \node_1.buffer_full_out , \node_1.receiving_data , 
        \node_1.sending_data , \node_1.data_in , \node_1.data_out  );
  input [15:0] \local_node.data_in ;
  output [15:0] \local_node.data_out ;
  input [15:0] \node_0.data_in ;
  output [15:0] \node_0.data_out ;
  input [15:0] \node_1.data_in ;
  output [15:0] \node_1.data_out ;
  input \clk.clk , \reset.reset , \local_node.buffer_full_in ,
         \local_node.receiving_data , \node_0.buffer_full_in ,
         \node_0.receiving_data , \node_1.buffer_full_in ,
         \node_1.receiving_data ;
  output \local_node.buffer_full_out , \local_node.sending_data ,
         \node_0.buffer_full_out , \node_0.sending_data ,
         \node_1.buffer_full_out , \node_1.sending_data ;
  inout \local_node.clk ,  \node_0.clk ,  \node_1.clk ;
  wire   \buffer_out[2][15] , \buffer_out[2][14] , \buffer_out[2][13] ,
         \buffer_out[2][12] , \buffer_out[2][11] , \buffer_out[2][10] ,
         \buffer_out[2][9] , \buffer_out[2][8] , \buffer_out[2][7] ,
         \buffer_out[2][6] , \buffer_out[2][5] , \buffer_out[2][4] ,
         \buffer_out[2][3] , \buffer_out[2][2] , \buffer_out[2][1] ,
         \buffer_out[2][0] , \buffer_out[1][15] , \buffer_out[1][14] ,
         \buffer_out[1][13] , \buffer_out[1][12] , \buffer_out[1][11] ,
         \buffer_out[1][10] , \buffer_out[1][9] , \buffer_out[1][8] ,
         \buffer_out[1][7] , \buffer_out[1][6] , \buffer_out[1][5] ,
         \buffer_out[1][4] , \buffer_out[1][3] , \buffer_out[1][2] ,
         \buffer_out[1][1] , \buffer_out[1][0] , \buffer_out[0][15] ,
         \buffer_out[0][14] , \buffer_out[0][13] , \buffer_out[0][12] ,
         \buffer_out[0][11] , \buffer_out[0][10] , \buffer_out[0][9] ,
         \buffer_out[0][8] , \buffer_out[0][7] , \buffer_out[0][6] ,
         \buffer_out[0][5] , \buffer_out[0][4] , \buffer_out[0][3] ,
         \buffer_out[0][2] , \buffer_out[0][1] , \buffer_out[0][0] ,
         \next_buffer_out[2][15] , \next_buffer_out[2][14] ,
         \next_buffer_out[2][13] , \next_buffer_out[2][12] ,
         \next_buffer_out[2][11] , \next_buffer_out[2][10] ,
         \next_buffer_out[2][9] , \next_buffer_out[2][8] ,
         \next_buffer_out[2][7] , \next_buffer_out[2][6] ,
         \next_buffer_out[2][5] , \next_buffer_out[2][4] ,
         \next_buffer_out[2][3] , \next_buffer_out[2][2] ,
         \next_buffer_out[2][1] , \next_buffer_out[2][0] ,
         \next_buffer_out[1][15] , \next_buffer_out[1][14] ,
         \next_buffer_out[1][13] , \next_buffer_out[1][12] ,
         \next_buffer_out[1][11] , \next_buffer_out[1][10] ,
         \next_buffer_out[1][9] , \next_buffer_out[1][8] ,
         \next_buffer_out[1][7] , \next_buffer_out[1][6] ,
         \next_buffer_out[1][5] , \next_buffer_out[1][4] ,
         \next_buffer_out[1][3] , \next_buffer_out[1][2] ,
         \next_buffer_out[1][1] , \next_buffer_out[1][0] ,
         \next_buffer_out[0][15] , \next_buffer_out[0][14] ,
         \next_buffer_out[0][13] , \next_buffer_out[0][12] ,
         \next_buffer_out[0][11] , \next_buffer_out[0][10] ,
         \next_buffer_out[0][9] , \next_buffer_out[0][8] ,
         \next_buffer_out[0][7] , \next_buffer_out[0][6] ,
         \next_buffer_out[0][5] , \next_buffer_out[0][4] ,
         \next_buffer_out[0][3] , \next_buffer_out[0][2] ,
         \next_buffer_out[0][1] , \next_buffer_out[0][0] ;
  wire   [2:0] buffer_full_in;
  wire   [2:0] receiving_data;
  wire   [2:0] pop_v;
  wire   [2:0] data_valid;
  wire   [2:0] next_data_valid;
  wire   [1:0] grant_1;
  wire   [1:0] grant_2;
  tri   \local_node.buffer_full_in ;
  tri   \local_node.buffer_full_out ;
  tri   \local_node.receiving_data ;
  tri   \local_node.sending_data ;
  tri   [15:0] \local_node.data_in ;
  tri   [15:0] \local_node.data_out ;

  converter_out_I_n_node_interface_dut_ c2 ( .\n.buffer_full_in (
        \local_node.buffer_full_in ), .\n.receiving_data (
        \local_node.receiving_data ), .\n.data_in (\local_node.data_in ), 
        .\n.buffer_full_out (\local_node.buffer_full_out ), .\n.sending_data (
        \local_node.sending_data ), .\n.data_out (\local_node.data_out ), 
        .buffer_full_in(1'b0), .receiving_data(1'b0), .data_in({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  fifo_kev_63 \genblk1[0].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[0]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[0]), .data_out({\buffer_out[0][15] , 
        \buffer_out[0][14] , \buffer_out[0][13] , \buffer_out[0][12] , 
        \buffer_out[0][11] , \buffer_out[0][10] , \buffer_out[0][9] , 
        \buffer_out[0][8] , \buffer_out[0][7] , \buffer_out[0][6] , 
        \buffer_out[0][5] , \buffer_out[0][4] , \buffer_out[0][3] , 
        \buffer_out[0][2] , \buffer_out[0][1] , \buffer_out[0][0] }), 
        .next_data_out({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] , 
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .next_data_valid(
        next_data_valid[0]) );
  address_counter_63 \genblk1[0].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] }), 
        .buffer_data_valid(next_data_valid[0]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .buffer_pop(
        pop_v[0]), .receiving_data(1'b0) );
  fifo_kev_62 \genblk1[1].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[1]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[1]), .data_out({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), 
        .next_data_out({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] , 
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .next_data_valid(
        next_data_valid[1]) );
  address_counter_62 \genblk1[1].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] }), 
        .buffer_data_valid(next_data_valid[1]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .buffer_pop(
        pop_v[1]), .receiving_data(1'b0) );
  fifo_kev_61 \genblk1[2].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[2]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[2]), .data_out({\buffer_out[2][15] , 
        \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] , 
        \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] , 
        \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] , 
        \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] , 
        \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] }), 
        .next_data_out({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] , 
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .next_data_valid(
        next_data_valid[2]) );
  address_counter_61 \genblk1[2].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] }), 
        .buffer_data_valid(next_data_valid[2]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .buffer_pop(
        pop_v[2]), .receiving_data(1'b0) );
  converter_out_I_n_node_interface_dut_ \genblk2.c0  ( .\n.buffer_full_in (
        \node_0.buffer_full_in ), .\n.receiving_data (\node_0.receiving_data ), 
        .\n.data_in (\node_0.data_in ), .\n.buffer_full_out (
        \node_0.buffer_full_out ), .\n.sending_data (\node_0.sending_data ), 
        .\n.data_out (\node_0.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_in_I_n_node_interface_dut__23 \genblk2.c1  ( .\n.buffer_full_in (
        \node_1.buffer_full_in ), .\n.receiving_data (\node_1.receiving_data ), 
        .\n.data_in (\node_1.data_in ), .\n.buffer_full_out (
        \node_1.buffer_full_out ), .\n.sending_data (\node_1.sending_data ), 
        .\n.data_out (\node_1.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  controller3_nw \genblk2.nw  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .packet_addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .local_addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .packet_valid(data_valid), .buffer_full_in({1'b0, 1'b0, 
        1'b0}), .grant_1(grant_1), .grant_2(grant_2), .pop_v(pop_v) );
  mux2_1_23 \genblk2.mux_w  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[2][15] , 
        \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] , 
        \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] , 
        \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] , 
        \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] , 
        \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] }), 
        .select0(grant_1[0]), .select1(grant_1[1]) );
  mux2_1_22 \genblk2.mux_l  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), 
        .select0(grant_2[0]), .select1(grant_2[1]) );
endmodule


module fifo_kev_60 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_121 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_60 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_121 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_120 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_60 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_120 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_60_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_60 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_60 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_60 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_60_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_59 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_119 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_59 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_119 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_118 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_59 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_118 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_59_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_59 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_59 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_59 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_59_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_58 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_117 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_58 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_117 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_116 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_58 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_116 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_58_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_58 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_58 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_58 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_58_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module flipflop_BITS2_21 ( clk, data_i, data_o );
  input [1:0] data_i;
  output [1:0] data_o;
  input clk;


  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS2_21 ( clk, enable_i, reset, data_i, data_o );
  input [1:0] data_i;
  input [1:0] data_o;
  input clk, enable_i, reset;
  wire   n10, n11, n1, n5, n7, n8, n9;
  wire   [1:0] write_data;

  AOI22X1 U5 ( .IN1(enable_i), .IN2(data_i[1]), .IN3(n10), .IN4(n1), .QN(n9)
         );
  AOI22X1 U6 ( .IN1(data_i[0]), .IN2(enable_i), .IN3(n11), .IN4(n1), .QN(n8)
         );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n9), .QN(write_data[1]) );
  NOR2X0 U4 ( .IN1(reset), .IN2(n8), .QN(write_data[0]) );
  AND2X1 U7 ( .IN1(data_o[1]), .IN2(n7), .Q(n10) );
  AND2X1 U8 ( .IN1(data_o[0]), .IN2(n5), .Q(n11) );
  flipflop_BITS2_21 FF ( .clk(clk), .data_i(write_data), .data_o({n7, n5}) );
endmodule


module flipflop_BITS1_85 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_85 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_85 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter2_21 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [1:0] request;
  output [1:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   tail_en, n1, n2;
  wire   [1:0] req_i;
  wire   [1:0] req_o;

  AND3X1 U10 ( .IN1(request[1]), .IN2(n1), .IN3(n2), .Q(grant[1]) );
  AND3X1 U11 ( .IN1(request[0]), .IN2(n2), .IN3(request[1]), .Q(tail_en) );
  INVX0 U6 ( .INP(request[0]), .ZN(n1) );
  NOR2X0 U7 ( .IN1(buffer_full_i), .IN2(n1), .QN(grant[0]) );
  INVX0 U8 ( .INP(buffer_full_i), .ZN(n2) );
  OA21X1 U9 ( .IN1(request[1]), .IN2(request[0]), .IN3(n2), .Q(grant_v_o) );
  register_BITS2_21 req_record ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i({1'b1, 1'b0}), .data_o({1'b0, 1'b0}) );
  register_BITS1_85 tail ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i(1'b1), .data_o(1'b0) );
endmodule


module flipflop_BITS2_20 ( clk, data_i, data_o );
  input [1:0] data_i;
  output [1:0] data_o;
  input clk;


  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS2_20 ( clk, enable_i, reset, data_i, data_o );
  input [1:0] data_i;
  input [1:0] data_o;
  input clk, enable_i, reset;
  wire   n10, n11, n1, n5, n7, n8, n9;
  wire   [1:0] write_data;

  AOI22X1 U5 ( .IN1(enable_i), .IN2(data_i[1]), .IN3(n10), .IN4(n1), .QN(n9)
         );
  AOI22X1 U6 ( .IN1(data_i[0]), .IN2(enable_i), .IN3(n11), .IN4(n1), .QN(n8)
         );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n9), .QN(write_data[1]) );
  NOR2X0 U4 ( .IN1(reset), .IN2(n8), .QN(write_data[0]) );
  AND2X1 U7 ( .IN1(data_o[1]), .IN2(n7), .Q(n10) );
  AND2X1 U8 ( .IN1(data_o[0]), .IN2(n5), .Q(n11) );
  flipflop_BITS2_20 FF ( .clk(clk), .data_i(write_data), .data_o({n7, n5}) );
endmodule


module flipflop_BITS1_84 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_84 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_84 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter2_20 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [1:0] request;
  output [1:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   tail_en, n1, n2;
  wire   [1:0] req_i;
  wire   [1:0] req_o;

  AND3X1 U10 ( .IN1(request[1]), .IN2(n1), .IN3(n2), .Q(grant[1]) );
  AND3X1 U11 ( .IN1(request[0]), .IN2(n2), .IN3(request[1]), .Q(tail_en) );
  INVX0 U6 ( .INP(request[0]), .ZN(n1) );
  NOR2X0 U7 ( .IN1(buffer_full_i), .IN2(n1), .QN(grant[0]) );
  INVX0 U8 ( .INP(buffer_full_i), .ZN(n2) );
  OA21X1 U9 ( .IN1(request[1]), .IN2(request[0]), .IN3(n2), .Q(grant_v_o) );
  register_BITS2_20 req_record ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i({1'b1, 1'b0}), .data_o({1'b0, 1'b0}) );
  register_BITS1_84 tail ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i(1'b1), .data_o(1'b0) );
endmodule


module dccl_60 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_59 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_58 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module controller3_ne ( clk, rst, .packet_addr({\packet_addr[2][7] , 
        \packet_addr[2][6] , \packet_addr[2][5] , \packet_addr[2][4] , 
        \packet_addr[2][3] , \packet_addr[2][2] , \packet_addr[2][1] , 
        \packet_addr[2][0] , \packet_addr[1][7] , \packet_addr[1][6] , 
        \packet_addr[1][5] , \packet_addr[1][4] , \packet_addr[1][3] , 
        \packet_addr[1][2] , \packet_addr[1][1] , \packet_addr[1][0] , 
        \packet_addr[0][7] , \packet_addr[0][6] , \packet_addr[0][5] , 
        \packet_addr[0][4] , \packet_addr[0][3] , \packet_addr[0][2] , 
        \packet_addr[0][1] , \packet_addr[0][0] }), local_addr, packet_valid, 
        buffer_full_in, grant_1, grant_2, grant_v, pop_v );
  input [7:0] local_addr;
  input [2:0] packet_valid;
  input [2:0] buffer_full_in;
  output [1:0] grant_1;
  output [1:0] grant_2;
  output [2:0] grant_v;
  output [2:0] pop_v;
  input clk, rst, \packet_addr[2][7] , \packet_addr[2][6] ,
         \packet_addr[2][5] , \packet_addr[2][4] , \packet_addr[2][3] ,
         \packet_addr[2][2] , \packet_addr[2][1] , \packet_addr[2][0] ,
         \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] ,
         \packet_addr[1][4] , \packet_addr[1][3] , \packet_addr[1][2] ,
         \packet_addr[1][1] , \packet_addr[1][0] , \packet_addr[0][7] ,
         \packet_addr[0][6] , \packet_addr[0][5] , \packet_addr[0][4] ,
         \packet_addr[0][3] , \packet_addr[0][2] , \packet_addr[0][1] ,
         \packet_addr[0][0] ;
  wire   \grant_2[1] , \request[2][1] , \request[2][0] , \request[1][1] ,
         \request[1][0] , \request[0][0] , n1;
  assign pop_v[1] = \grant_2[1] ;
  assign grant_2[1] = \grant_2[1] ;

  OR2X1 U3 ( .IN1(grant_v[0]), .IN2(grant_1[1]), .Q(pop_v[2]) );
  OR2X1 U4 ( .IN1(grant_1[0]), .IN2(grant_2[0]), .Q(pop_v[0]) );
  NOR2X0 U1 ( .IN1(n1), .IN2(buffer_full_in[0]), .QN(grant_v[0]) );
  INVX0 U2 ( .INP(\request[0][0] ), .ZN(n1) );
  arbiter2_21 arbiter_w ( .clk(clk), .rst(rst), .request({\request[1][1] , 
        \request[1][0] }), .buffer_full_i(buffer_full_in[1]), .grant(grant_1), 
        .grant_v_o(grant_v[1]) );
  arbiter2_20 arbiter_l ( .clk(clk), .rst(rst), .request({\request[2][1] , 
        \request[2][0] }), .buffer_full_i(buffer_full_in[2]), .grant({
        \grant_2[1] , grant_2[0]}), .grant_v_o(grant_v[2]) );
  dccl_60 dccl_s ( .packet_addr_y_i({\packet_addr[0][3] , \packet_addr[0][2] , 
        \packet_addr[0][1] , \packet_addr[0][0] }), .packet_addr_x_i({
        \packet_addr[0][7] , \packet_addr[0][6] , \packet_addr[0][5] , 
        \packet_addr[0][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[0]), 
        .west_req(\request[1][0] ), .local_req(\request[2][0] ) );
  dccl_59 dccl_w ( .packet_addr_y_i({\packet_addr[1][3] , \packet_addr[1][2] , 
        \packet_addr[1][1] , \packet_addr[1][0] }), .packet_addr_x_i({
        \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] , 
        \packet_addr[1][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[1]), 
        .local_req(\request[2][1] ) );
  dccl_58 dccl_l ( .packet_addr_y_i({\packet_addr[2][3] , \packet_addr[2][2] , 
        \packet_addr[2][1] , \packet_addr[2][0] }), .packet_addr_x_i({
        \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] , 
        \packet_addr[2][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[2]), 
        .south_req(\request[0][0] ), .west_req(\request[1][1] ) );
endmodule


module mux2_1_21 ( data0, data1, select0, select1, data_o );
  input [15:0] data0;
  input [15:0] data1;
  output [15:0] data_o;
  input select0, select1;
  wire   n1, n4, n5;

  AO22X1 U4 ( .IN1(data1[9]), .IN2(n5), .IN3(data0[9]), .IN4(n4), .Q(data_o[9]) );
  AO22X1 U5 ( .IN1(data1[8]), .IN2(n5), .IN3(data0[8]), .IN4(n4), .Q(data_o[8]) );
  AO22X1 U6 ( .IN1(data1[7]), .IN2(n5), .IN3(data0[7]), .IN4(n4), .Q(data_o[7]) );
  AO22X1 U7 ( .IN1(data1[6]), .IN2(n5), .IN3(data0[6]), .IN4(n4), .Q(data_o[6]) );
  AO22X1 U8 ( .IN1(data1[5]), .IN2(n5), .IN3(data0[5]), .IN4(n4), .Q(data_o[5]) );
  AO22X1 U9 ( .IN1(data1[4]), .IN2(n5), .IN3(data0[4]), .IN4(n4), .Q(data_o[4]) );
  AO22X1 U10 ( .IN1(data1[3]), .IN2(n5), .IN3(data0[3]), .IN4(n4), .Q(
        data_o[3]) );
  AO22X1 U11 ( .IN1(data1[2]), .IN2(n5), .IN3(data0[2]), .IN4(n4), .Q(
        data_o[2]) );
  AO22X1 U12 ( .IN1(data1[1]), .IN2(n5), .IN3(data0[1]), .IN4(n4), .Q(
        data_o[1]) );
  AO22X1 U13 ( .IN1(data1[15]), .IN2(n5), .IN3(data0[15]), .IN4(n4), .Q(
        data_o[15]) );
  AO22X1 U14 ( .IN1(data1[14]), .IN2(n5), .IN3(data0[14]), .IN4(n4), .Q(
        data_o[14]) );
  AO22X1 U15 ( .IN1(data1[13]), .IN2(n5), .IN3(data0[13]), .IN4(n4), .Q(
        data_o[13]) );
  AO22X1 U16 ( .IN1(data1[12]), .IN2(n5), .IN3(data0[12]), .IN4(n4), .Q(
        data_o[12]) );
  AO22X1 U17 ( .IN1(data1[11]), .IN2(n5), .IN3(data0[11]), .IN4(n4), .Q(
        data_o[11]) );
  AO22X1 U18 ( .IN1(data1[10]), .IN2(n5), .IN3(data0[10]), .IN4(n4), .Q(
        data_o[10]) );
  AO22X1 U19 ( .IN1(data1[0]), .IN2(n5), .IN3(data0[0]), .IN4(n4), .Q(
        data_o[0]) );
  INVX0 U2 ( .INP(select1), .ZN(n1) );
  AND2X1 U3 ( .IN1(select0), .IN2(n1), .Q(n4) );
  NOR2X0 U20 ( .IN1(n1), .IN2(select0), .QN(n5) );
endmodule


module mux2_1_20 ( data0, data1, select0, select1, data_o );
  input [15:0] data0;
  input [15:0] data1;
  output [15:0] data_o;
  input select0, select1;
  wire   n1, n4, n5;

  AO22X1 U4 ( .IN1(data1[9]), .IN2(n5), .IN3(data0[9]), .IN4(n4), .Q(data_o[9]) );
  AO22X1 U5 ( .IN1(data1[8]), .IN2(n5), .IN3(data0[8]), .IN4(n4), .Q(data_o[8]) );
  AO22X1 U6 ( .IN1(data1[7]), .IN2(n5), .IN3(data0[7]), .IN4(n4), .Q(data_o[7]) );
  AO22X1 U7 ( .IN1(data1[6]), .IN2(n5), .IN3(data0[6]), .IN4(n4), .Q(data_o[6]) );
  AO22X1 U8 ( .IN1(data1[5]), .IN2(n5), .IN3(data0[5]), .IN4(n4), .Q(data_o[5]) );
  AO22X1 U9 ( .IN1(data1[4]), .IN2(n5), .IN3(data0[4]), .IN4(n4), .Q(data_o[4]) );
  AO22X1 U10 ( .IN1(data1[3]), .IN2(n5), .IN3(data0[3]), .IN4(n4), .Q(
        data_o[3]) );
  AO22X1 U11 ( .IN1(data1[2]), .IN2(n5), .IN3(data0[2]), .IN4(n4), .Q(
        data_o[2]) );
  AO22X1 U12 ( .IN1(data1[1]), .IN2(n5), .IN3(data0[1]), .IN4(n4), .Q(
        data_o[1]) );
  AO22X1 U13 ( .IN1(data1[15]), .IN2(n5), .IN3(data0[15]), .IN4(n4), .Q(
        data_o[15]) );
  AO22X1 U14 ( .IN1(data1[14]), .IN2(n5), .IN3(data0[14]), .IN4(n4), .Q(
        data_o[14]) );
  AO22X1 U15 ( .IN1(data1[13]), .IN2(n5), .IN3(data0[13]), .IN4(n4), .Q(
        data_o[13]) );
  AO22X1 U16 ( .IN1(data1[12]), .IN2(n5), .IN3(data0[12]), .IN4(n4), .Q(
        data_o[12]) );
  AO22X1 U17 ( .IN1(data1[11]), .IN2(n5), .IN3(data0[11]), .IN4(n4), .Q(
        data_o[11]) );
  AO22X1 U18 ( .IN1(data1[10]), .IN2(n5), .IN3(data0[10]), .IN4(n4), .Q(
        data_o[10]) );
  AO22X1 U19 ( .IN1(data1[0]), .IN2(n5), .IN3(data0[0]), .IN4(n4), .Q(
        data_o[0]) );
  INVX0 U2 ( .INP(select1), .ZN(n1) );
  AND2X1 U3 ( .IN1(select0), .IN2(n1), .Q(n4) );
  NOR2X0 U20 ( .IN1(n1), .IN2(select0), .QN(n5) );
endmodule



    module node3_NODE_X3_NODE_Y0I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__ ( 
        \clk.clk , \reset.reset , \local_node.clk , 
        \local_node.buffer_full_in , \local_node.buffer_full_out , 
        \local_node.receiving_data , \local_node.sending_data , 
        \local_node.data_in , \local_node.data_out , \node_0.clk , 
        \node_0.buffer_full_in , \node_0.buffer_full_out , 
        \node_0.receiving_data , \node_0.sending_data , \node_0.data_in , 
        \node_0.data_out , \node_1.clk , \node_1.buffer_full_in , 
        \node_1.buffer_full_out , \node_1.receiving_data , 
        \node_1.sending_data , \node_1.data_in , \node_1.data_out  );
  input [15:0] \local_node.data_in ;
  output [15:0] \local_node.data_out ;
  input [15:0] \node_0.data_in ;
  output [15:0] \node_0.data_out ;
  input [15:0] \node_1.data_in ;
  output [15:0] \node_1.data_out ;
  input \clk.clk , \reset.reset , \local_node.buffer_full_in ,
         \local_node.receiving_data , \node_0.buffer_full_in ,
         \node_0.receiving_data , \node_1.buffer_full_in ,
         \node_1.receiving_data ;
  output \local_node.buffer_full_out , \local_node.sending_data ,
         \node_0.buffer_full_out , \node_0.sending_data ,
         \node_1.buffer_full_out , \node_1.sending_data ;
  inout \local_node.clk ,  \node_0.clk ,  \node_1.clk ;
  wire   \buffer_out[2][15] , \buffer_out[2][14] , \buffer_out[2][13] ,
         \buffer_out[2][12] , \buffer_out[2][11] , \buffer_out[2][10] ,
         \buffer_out[2][9] , \buffer_out[2][8] , \buffer_out[2][7] ,
         \buffer_out[2][6] , \buffer_out[2][5] , \buffer_out[2][4] ,
         \buffer_out[2][3] , \buffer_out[2][2] , \buffer_out[2][1] ,
         \buffer_out[2][0] , \buffer_out[1][15] , \buffer_out[1][14] ,
         \buffer_out[1][13] , \buffer_out[1][12] , \buffer_out[1][11] ,
         \buffer_out[1][10] , \buffer_out[1][9] , \buffer_out[1][8] ,
         \buffer_out[1][7] , \buffer_out[1][6] , \buffer_out[1][5] ,
         \buffer_out[1][4] , \buffer_out[1][3] , \buffer_out[1][2] ,
         \buffer_out[1][1] , \buffer_out[1][0] , \buffer_out[0][15] ,
         \buffer_out[0][14] , \buffer_out[0][13] , \buffer_out[0][12] ,
         \buffer_out[0][11] , \buffer_out[0][10] , \buffer_out[0][9] ,
         \buffer_out[0][8] , \buffer_out[0][7] , \buffer_out[0][6] ,
         \buffer_out[0][5] , \buffer_out[0][4] , \buffer_out[0][3] ,
         \buffer_out[0][2] , \buffer_out[0][1] , \buffer_out[0][0] ,
         \next_buffer_out[2][15] , \next_buffer_out[2][14] ,
         \next_buffer_out[2][13] , \next_buffer_out[2][12] ,
         \next_buffer_out[2][11] , \next_buffer_out[2][10] ,
         \next_buffer_out[2][9] , \next_buffer_out[2][8] ,
         \next_buffer_out[2][7] , \next_buffer_out[2][6] ,
         \next_buffer_out[2][5] , \next_buffer_out[2][4] ,
         \next_buffer_out[2][3] , \next_buffer_out[2][2] ,
         \next_buffer_out[2][1] , \next_buffer_out[2][0] ,
         \next_buffer_out[1][15] , \next_buffer_out[1][14] ,
         \next_buffer_out[1][13] , \next_buffer_out[1][12] ,
         \next_buffer_out[1][11] , \next_buffer_out[1][10] ,
         \next_buffer_out[1][9] , \next_buffer_out[1][8] ,
         \next_buffer_out[1][7] , \next_buffer_out[1][6] ,
         \next_buffer_out[1][5] , \next_buffer_out[1][4] ,
         \next_buffer_out[1][3] , \next_buffer_out[1][2] ,
         \next_buffer_out[1][1] , \next_buffer_out[1][0] ,
         \next_buffer_out[0][15] , \next_buffer_out[0][14] ,
         \next_buffer_out[0][13] , \next_buffer_out[0][12] ,
         \next_buffer_out[0][11] , \next_buffer_out[0][10] ,
         \next_buffer_out[0][9] , \next_buffer_out[0][8] ,
         \next_buffer_out[0][7] , \next_buffer_out[0][6] ,
         \next_buffer_out[0][5] , \next_buffer_out[0][4] ,
         \next_buffer_out[0][3] , \next_buffer_out[0][2] ,
         \next_buffer_out[0][1] , \next_buffer_out[0][0] ;
  wire   [2:0] buffer_full_in;
  wire   [2:0] receiving_data;
  wire   [2:0] pop_v;
  wire   [2:0] data_valid;
  wire   [2:0] next_data_valid;
  wire   [1:0] grant_1;
  wire   [1:0] grant_2;
  tri   \local_node.buffer_full_in ;
  tri   \local_node.buffer_full_out ;
  tri   \local_node.receiving_data ;
  tri   \local_node.sending_data ;
  tri   [15:0] \local_node.data_in ;
  tri   [15:0] \local_node.data_out ;

  converter_out_I_n_node_interface_dut_ c2 ( .\n.buffer_full_in (
        \local_node.buffer_full_in ), .\n.receiving_data (
        \local_node.receiving_data ), .\n.data_in (\local_node.data_in ), 
        .\n.buffer_full_out (\local_node.buffer_full_out ), .\n.sending_data (
        \local_node.sending_data ), .\n.data_out (\local_node.data_out ), 
        .buffer_full_in(1'b0), .receiving_data(1'b0), .data_in({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  fifo_kev_60 \genblk1[0].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[0]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[0]), .data_out({\buffer_out[0][15] , 
        \buffer_out[0][14] , \buffer_out[0][13] , \buffer_out[0][12] , 
        \buffer_out[0][11] , \buffer_out[0][10] , \buffer_out[0][9] , 
        \buffer_out[0][8] , \buffer_out[0][7] , \buffer_out[0][6] , 
        \buffer_out[0][5] , \buffer_out[0][4] , \buffer_out[0][3] , 
        \buffer_out[0][2] , \buffer_out[0][1] , \buffer_out[0][0] }), 
        .next_data_out({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] , 
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .next_data_valid(
        next_data_valid[0]) );
  address_counter_60 \genblk1[0].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] }), 
        .buffer_data_valid(next_data_valid[0]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .buffer_pop(
        pop_v[0]), .receiving_data(1'b0) );
  fifo_kev_59 \genblk1[1].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[1]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[1]), .data_out({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), 
        .next_data_out({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] , 
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .next_data_valid(
        next_data_valid[1]) );
  address_counter_59 \genblk1[1].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] }), 
        .buffer_data_valid(next_data_valid[1]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .buffer_pop(
        pop_v[1]), .receiving_data(1'b0) );
  fifo_kev_58 \genblk1[2].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[2]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[2]), .data_out({\buffer_out[2][15] , 
        \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] , 
        \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] , 
        \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] , 
        \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] , 
        \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] }), 
        .next_data_out({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] , 
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .next_data_valid(
        next_data_valid[2]) );
  address_counter_58 \genblk1[2].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] }), 
        .buffer_data_valid(next_data_valid[2]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .buffer_pop(
        pop_v[2]), .receiving_data(1'b0) );
  converter_out_I_n_node_interface_dut_ \genblk2.c0  ( .\n.buffer_full_in (
        \node_0.buffer_full_in ), .\n.receiving_data (\node_0.receiving_data ), 
        .\n.data_in (\node_0.data_in ), .\n.buffer_full_out (
        \node_0.buffer_full_out ), .\n.sending_data (\node_0.sending_data ), 
        .\n.data_out (\node_0.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_out_I_n_node_interface_dut_ \genblk2.c1  ( .\n.buffer_full_in (
        \node_1.buffer_full_in ), .\n.receiving_data (\node_1.receiving_data ), 
        .\n.data_in (\node_1.data_in ), .\n.buffer_full_out (
        \node_1.buffer_full_out ), .\n.sending_data (\node_1.sending_data ), 
        .\n.data_out (\node_1.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  controller3_ne \genblk2.ne  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .packet_addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .local_addr({1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 
        1'b0, 1'b0}), .packet_valid(data_valid), .buffer_full_in({1'b0, 1'b0, 
        1'b0}), .grant_1(grant_1), .grant_2(grant_2), .pop_v(pop_v) );
  mux2_1_21 \genblk2.mux_e  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[2][15] , 
        \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] , 
        \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] , 
        \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] , 
        \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] , 
        \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] }), 
        .select0(grant_1[0]), .select1(grant_1[1]) );
  mux2_1_20 \genblk2.mux_l  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), 
        .select0(grant_2[0]), .select1(grant_2[1]) );
endmodule


module fifo_kev_57 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_115 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_57 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_115 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_114 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_57 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_114 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_57_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_57 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_57 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_57 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_57_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_56 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_113 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_56 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_113 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_112 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_56 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_112 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_56_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_56 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_56 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_56 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_56_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_55 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_111 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_55 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_111 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_110 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_55 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_110 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_55_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_55 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_55 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_55 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_55_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module converter_in_I_n_node_interface_dut__22 ( \n.buffer_full_in , 
        \n.receiving_data , \n.data_in , \n.buffer_full_out , \n.sending_data , 
        \n.data_out , buffer_full_out, sending_data, data_out, buffer_full_in, 
        receiving_data, data_in );
  input [15:0] \n.data_in ;
  output [15:0] \n.data_out ;
  output [15:0] data_out;
  input [15:0] data_in;
  input \n.buffer_full_in , \n.receiving_data , buffer_full_in, receiving_data;
  output \n.buffer_full_out , \n.sending_data , buffer_full_out, sending_data;
  wire   \n.buffer_full_in , \n.receiving_data , buffer_full_in,
         receiving_data;
  assign buffer_full_out = \n.buffer_full_in ;
  assign sending_data = \n.receiving_data ;
  assign data_out[15] = \n.data_in  [15];
  assign data_out[14] = \n.data_in  [14];
  assign data_out[13] = \n.data_in  [13];
  assign data_out[12] = \n.data_in  [12];
  assign data_out[11] = \n.data_in  [11];
  assign data_out[10] = \n.data_in  [10];
  assign data_out[9] = \n.data_in  [9];
  assign data_out[8] = \n.data_in  [8];
  assign data_out[7] = \n.data_in  [7];
  assign data_out[6] = \n.data_in  [6];
  assign data_out[5] = \n.data_in  [5];
  assign data_out[4] = \n.data_in  [4];
  assign data_out[3] = \n.data_in  [3];
  assign data_out[2] = \n.data_in  [2];
  assign data_out[1] = \n.data_in  [1];
  assign data_out[0] = \n.data_in  [0];
  assign \n.buffer_full_out  = buffer_full_in;
  assign \n.sending_data  = receiving_data;
  assign \n.data_out  [15] = data_in[15];
  assign \n.data_out  [14] = data_in[14];
  assign \n.data_out  [13] = data_in[13];
  assign \n.data_out  [12] = data_in[12];
  assign \n.data_out  [11] = data_in[11];
  assign \n.data_out  [10] = data_in[10];
  assign \n.data_out  [9] = data_in[9];
  assign \n.data_out  [8] = data_in[8];
  assign \n.data_out  [7] = data_in[7];
  assign \n.data_out  [6] = data_in[6];
  assign \n.data_out  [5] = data_in[5];
  assign \n.data_out  [4] = data_in[4];
  assign \n.data_out  [3] = data_in[3];
  assign \n.data_out  [2] = data_in[2];
  assign \n.data_out  [1] = data_in[1];
  assign \n.data_out  [0] = data_in[0];

endmodule


module converter_in_I_n_node_interface_dut__21 ( \n.buffer_full_in , 
        \n.receiving_data , \n.data_in , \n.buffer_full_out , \n.sending_data , 
        \n.data_out , buffer_full_out, sending_data, data_out, buffer_full_in, 
        receiving_data, data_in );
  input [15:0] \n.data_in ;
  output [15:0] \n.data_out ;
  output [15:0] data_out;
  input [15:0] data_in;
  input \n.buffer_full_in , \n.receiving_data , buffer_full_in, receiving_data;
  output \n.buffer_full_out , \n.sending_data , buffer_full_out, sending_data;
  wire   \n.buffer_full_in , \n.receiving_data , buffer_full_in,
         receiving_data;
  assign buffer_full_out = \n.buffer_full_in ;
  assign sending_data = \n.receiving_data ;
  assign data_out[15] = \n.data_in  [15];
  assign data_out[14] = \n.data_in  [14];
  assign data_out[13] = \n.data_in  [13];
  assign data_out[12] = \n.data_in  [12];
  assign data_out[11] = \n.data_in  [11];
  assign data_out[10] = \n.data_in  [10];
  assign data_out[9] = \n.data_in  [9];
  assign data_out[8] = \n.data_in  [8];
  assign data_out[7] = \n.data_in  [7];
  assign data_out[6] = \n.data_in  [6];
  assign data_out[5] = \n.data_in  [5];
  assign data_out[4] = \n.data_in  [4];
  assign data_out[3] = \n.data_in  [3];
  assign data_out[2] = \n.data_in  [2];
  assign data_out[1] = \n.data_in  [1];
  assign data_out[0] = \n.data_in  [0];
  assign \n.buffer_full_out  = buffer_full_in;
  assign \n.sending_data  = receiving_data;
  assign \n.data_out  [15] = data_in[15];
  assign \n.data_out  [14] = data_in[14];
  assign \n.data_out  [13] = data_in[13];
  assign \n.data_out  [12] = data_in[12];
  assign \n.data_out  [11] = data_in[11];
  assign \n.data_out  [10] = data_in[10];
  assign \n.data_out  [9] = data_in[9];
  assign \n.data_out  [8] = data_in[8];
  assign \n.data_out  [7] = data_in[7];
  assign \n.data_out  [6] = data_in[6];
  assign \n.data_out  [5] = data_in[5];
  assign \n.data_out  [4] = data_in[4];
  assign \n.data_out  [3] = data_in[3];
  assign \n.data_out  [2] = data_in[2];
  assign \n.data_out  [1] = data_in[1];
  assign \n.data_out  [0] = data_in[0];

endmodule


module flipflop_BITS2_19 ( clk, data_i, data_o );
  input [1:0] data_i;
  output [1:0] data_o;
  input clk;


  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS2_19 ( clk, enable_i, reset, data_i, data_o );
  input [1:0] data_i;
  input [1:0] data_o;
  input clk, enable_i, reset;
  wire   n10, n11, n1, n5, n7, n8, n9;
  wire   [1:0] write_data;

  AOI22X1 U5 ( .IN1(enable_i), .IN2(data_i[1]), .IN3(n10), .IN4(n1), .QN(n9)
         );
  AOI22X1 U6 ( .IN1(data_i[0]), .IN2(enable_i), .IN3(n11), .IN4(n1), .QN(n8)
         );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n9), .QN(write_data[1]) );
  NOR2X0 U4 ( .IN1(reset), .IN2(n8), .QN(write_data[0]) );
  AND2X1 U7 ( .IN1(data_o[1]), .IN2(n7), .Q(n10) );
  AND2X1 U8 ( .IN1(data_o[0]), .IN2(n5), .Q(n11) );
  flipflop_BITS2_19 FF ( .clk(clk), .data_i(write_data), .data_o({n7, n5}) );
endmodule


module flipflop_BITS1_83 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_83 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_83 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter2_19 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [1:0] request;
  output [1:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   tail_en, n1, n2;
  wire   [1:0] req_i;
  wire   [1:0] req_o;

  AND3X1 U10 ( .IN1(request[1]), .IN2(n1), .IN3(n2), .Q(grant[1]) );
  AND3X1 U11 ( .IN1(request[0]), .IN2(n2), .IN3(request[1]), .Q(tail_en) );
  INVX0 U6 ( .INP(request[0]), .ZN(n1) );
  NOR2X0 U7 ( .IN1(buffer_full_i), .IN2(n1), .QN(grant[0]) );
  INVX0 U8 ( .INP(buffer_full_i), .ZN(n2) );
  OA21X1 U9 ( .IN1(request[1]), .IN2(request[0]), .IN3(n2), .Q(grant_v_o) );
  register_BITS2_19 req_record ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i({1'b1, 1'b0}), .data_o({1'b0, 1'b0}) );
  register_BITS1_83 tail ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i(1'b1), .data_o(1'b0) );
endmodule


module flipflop_BITS2_18 ( clk, data_i, data_o );
  input [1:0] data_i;
  output [1:0] data_o;
  input clk;


  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS2_18 ( clk, enable_i, reset, data_i, data_o );
  input [1:0] data_i;
  input [1:0] data_o;
  input clk, enable_i, reset;
  wire   n10, n11, n1, n5, n7, n8, n9;
  wire   [1:0] write_data;

  AOI22X1 U5 ( .IN1(enable_i), .IN2(data_i[1]), .IN3(n10), .IN4(n1), .QN(n9)
         );
  AOI22X1 U6 ( .IN1(data_i[0]), .IN2(enable_i), .IN3(n11), .IN4(n1), .QN(n8)
         );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n9), .QN(write_data[1]) );
  NOR2X0 U4 ( .IN1(reset), .IN2(n8), .QN(write_data[0]) );
  AND2X1 U7 ( .IN1(data_o[1]), .IN2(n7), .Q(n10) );
  AND2X1 U8 ( .IN1(data_o[0]), .IN2(n5), .Q(n11) );
  flipflop_BITS2_18 FF ( .clk(clk), .data_i(write_data), .data_o({n7, n5}) );
endmodule


module flipflop_BITS1_82 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_82 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_82 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter2_18 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [1:0] request;
  output [1:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   tail_en, n1, n2;
  wire   [1:0] req_i;
  wire   [1:0] req_o;

  AND3X1 U10 ( .IN1(request[1]), .IN2(n1), .IN3(n2), .Q(grant[1]) );
  AND3X1 U11 ( .IN1(request[0]), .IN2(n2), .IN3(request[1]), .Q(tail_en) );
  INVX0 U6 ( .INP(request[0]), .ZN(n1) );
  NOR2X0 U7 ( .IN1(buffer_full_i), .IN2(n1), .QN(grant[0]) );
  INVX0 U8 ( .INP(buffer_full_i), .ZN(n2) );
  OA21X1 U9 ( .IN1(request[1]), .IN2(request[0]), .IN3(n2), .Q(grant_v_o) );
  register_BITS2_18 req_record ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i({1'b1, 1'b0}), .data_o({1'b0, 1'b0}) );
  register_BITS1_82 tail ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i(1'b1), .data_o(1'b0) );
endmodule


module dccl_57 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_56 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_55 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module controller3_sw ( clk, rst, .packet_addr({\packet_addr[2][7] , 
        \packet_addr[2][6] , \packet_addr[2][5] , \packet_addr[2][4] , 
        \packet_addr[2][3] , \packet_addr[2][2] , \packet_addr[2][1] , 
        \packet_addr[2][0] , \packet_addr[1][7] , \packet_addr[1][6] , 
        \packet_addr[1][5] , \packet_addr[1][4] , \packet_addr[1][3] , 
        \packet_addr[1][2] , \packet_addr[1][1] , \packet_addr[1][0] , 
        \packet_addr[0][7] , \packet_addr[0][6] , \packet_addr[0][5] , 
        \packet_addr[0][4] , \packet_addr[0][3] , \packet_addr[0][2] , 
        \packet_addr[0][1] , \packet_addr[0][0] }), local_addr, packet_valid, 
        buffer_full_in, grant_1, grant_2, grant_v, pop_v );
  input [7:0] local_addr;
  input [2:0] packet_valid;
  input [2:0] buffer_full_in;
  output [1:0] grant_1;
  output [1:0] grant_2;
  output [2:0] grant_v;
  output [2:0] pop_v;
  input clk, rst, \packet_addr[2][7] , \packet_addr[2][6] ,
         \packet_addr[2][5] , \packet_addr[2][4] , \packet_addr[2][3] ,
         \packet_addr[2][2] , \packet_addr[2][1] , \packet_addr[2][0] ,
         \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] ,
         \packet_addr[1][4] , \packet_addr[1][3] , \packet_addr[1][2] ,
         \packet_addr[1][1] , \packet_addr[1][0] , \packet_addr[0][7] ,
         \packet_addr[0][6] , \packet_addr[0][5] , \packet_addr[0][4] ,
         \packet_addr[0][3] , \packet_addr[0][2] , \packet_addr[0][1] ,
         \packet_addr[0][0] ;
  wire   \grant_2[1] , \request[2][1] , \request[2][0] , \request[1][1] ,
         \request[1][0] , \request[0][0] , n1;
  assign pop_v[1] = \grant_2[1] ;
  assign grant_2[1] = \grant_2[1] ;

  OR2X1 U3 ( .IN1(grant_v[0]), .IN2(grant_1[1]), .Q(pop_v[2]) );
  OR2X1 U4 ( .IN1(grant_1[0]), .IN2(grant_2[0]), .Q(pop_v[0]) );
  NOR2X0 U1 ( .IN1(n1), .IN2(buffer_full_in[0]), .QN(grant_v[0]) );
  INVX0 U2 ( .INP(\request[0][0] ), .ZN(n1) );
  arbiter2_19 arbiter_e ( .clk(clk), .rst(rst), .request({\request[1][1] , 
        \request[1][0] }), .buffer_full_i(buffer_full_in[1]), .grant(grant_1), 
        .grant_v_o(grant_v[1]) );
  arbiter2_18 arbiter_l ( .clk(clk), .rst(rst), .request({\request[2][1] , 
        \request[2][0] }), .buffer_full_i(buffer_full_in[2]), .grant({
        \grant_2[1] , grant_2[0]}), .grant_v_o(grant_v[2]) );
  dccl_57 dccl_n ( .packet_addr_y_i({\packet_addr[0][3] , \packet_addr[0][2] , 
        \packet_addr[0][1] , \packet_addr[0][0] }), .packet_addr_x_i({
        \packet_addr[0][7] , \packet_addr[0][6] , \packet_addr[0][5] , 
        \packet_addr[0][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[0]), 
        .east_req(\request[1][0] ), .local_req(\request[2][0] ) );
  dccl_56 dccl_e ( .packet_addr_y_i({\packet_addr[1][3] , \packet_addr[1][2] , 
        \packet_addr[1][1] , \packet_addr[1][0] }), .packet_addr_x_i({
        \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] , 
        \packet_addr[1][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[1]), 
        .local_req(\request[2][1] ) );
  dccl_55 dccl_l ( .packet_addr_y_i({\packet_addr[2][3] , \packet_addr[2][2] , 
        \packet_addr[2][1] , \packet_addr[2][0] }), .packet_addr_x_i({
        \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] , 
        \packet_addr[2][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[2]), 
        .north_req(\request[0][0] ), .east_req(\request[1][1] ) );
endmodule


module mux2_1_19 ( data0, data1, select0, select1, data_o );
  input [15:0] data0;
  input [15:0] data1;
  output [15:0] data_o;
  input select0, select1;
  wire   n1, n4, n5;

  AO22X1 U4 ( .IN1(data1[9]), .IN2(n5), .IN3(data0[9]), .IN4(n4), .Q(data_o[9]) );
  AO22X1 U5 ( .IN1(data1[8]), .IN2(n5), .IN3(data0[8]), .IN4(n4), .Q(data_o[8]) );
  AO22X1 U6 ( .IN1(data1[7]), .IN2(n5), .IN3(data0[7]), .IN4(n4), .Q(data_o[7]) );
  AO22X1 U7 ( .IN1(data1[6]), .IN2(n5), .IN3(data0[6]), .IN4(n4), .Q(data_o[6]) );
  AO22X1 U8 ( .IN1(data1[5]), .IN2(n5), .IN3(data0[5]), .IN4(n4), .Q(data_o[5]) );
  AO22X1 U9 ( .IN1(data1[4]), .IN2(n5), .IN3(data0[4]), .IN4(n4), .Q(data_o[4]) );
  AO22X1 U10 ( .IN1(data1[3]), .IN2(n5), .IN3(data0[3]), .IN4(n4), .Q(
        data_o[3]) );
  AO22X1 U11 ( .IN1(data1[2]), .IN2(n5), .IN3(data0[2]), .IN4(n4), .Q(
        data_o[2]) );
  AO22X1 U12 ( .IN1(data1[1]), .IN2(n5), .IN3(data0[1]), .IN4(n4), .Q(
        data_o[1]) );
  AO22X1 U13 ( .IN1(data1[15]), .IN2(n5), .IN3(data0[15]), .IN4(n4), .Q(
        data_o[15]) );
  AO22X1 U14 ( .IN1(data1[14]), .IN2(n5), .IN3(data0[14]), .IN4(n4), .Q(
        data_o[14]) );
  AO22X1 U15 ( .IN1(data1[13]), .IN2(n5), .IN3(data0[13]), .IN4(n4), .Q(
        data_o[13]) );
  AO22X1 U16 ( .IN1(data1[12]), .IN2(n5), .IN3(data0[12]), .IN4(n4), .Q(
        data_o[12]) );
  AO22X1 U17 ( .IN1(data1[11]), .IN2(n5), .IN3(data0[11]), .IN4(n4), .Q(
        data_o[11]) );
  AO22X1 U18 ( .IN1(data1[10]), .IN2(n5), .IN3(data0[10]), .IN4(n4), .Q(
        data_o[10]) );
  AO22X1 U19 ( .IN1(data1[0]), .IN2(n5), .IN3(data0[0]), .IN4(n4), .Q(
        data_o[0]) );
  INVX0 U2 ( .INP(select1), .ZN(n1) );
  AND2X1 U3 ( .IN1(select0), .IN2(n1), .Q(n4) );
  NOR2X0 U20 ( .IN1(n1), .IN2(select0), .QN(n5) );
endmodule


module mux2_1_18 ( data0, data1, select0, select1, data_o );
  input [15:0] data0;
  input [15:0] data1;
  output [15:0] data_o;
  input select0, select1;
  wire   n1, n4, n5;

  AO22X1 U4 ( .IN1(data1[9]), .IN2(n5), .IN3(data0[9]), .IN4(n4), .Q(data_o[9]) );
  AO22X1 U5 ( .IN1(data1[8]), .IN2(n5), .IN3(data0[8]), .IN4(n4), .Q(data_o[8]) );
  AO22X1 U6 ( .IN1(data1[7]), .IN2(n5), .IN3(data0[7]), .IN4(n4), .Q(data_o[7]) );
  AO22X1 U7 ( .IN1(data1[6]), .IN2(n5), .IN3(data0[6]), .IN4(n4), .Q(data_o[6]) );
  AO22X1 U8 ( .IN1(data1[5]), .IN2(n5), .IN3(data0[5]), .IN4(n4), .Q(data_o[5]) );
  AO22X1 U9 ( .IN1(data1[4]), .IN2(n5), .IN3(data0[4]), .IN4(n4), .Q(data_o[4]) );
  AO22X1 U10 ( .IN1(data1[3]), .IN2(n5), .IN3(data0[3]), .IN4(n4), .Q(
        data_o[3]) );
  AO22X1 U11 ( .IN1(data1[2]), .IN2(n5), .IN3(data0[2]), .IN4(n4), .Q(
        data_o[2]) );
  AO22X1 U12 ( .IN1(data1[1]), .IN2(n5), .IN3(data0[1]), .IN4(n4), .Q(
        data_o[1]) );
  AO22X1 U13 ( .IN1(data1[15]), .IN2(n5), .IN3(data0[15]), .IN4(n4), .Q(
        data_o[15]) );
  AO22X1 U14 ( .IN1(data1[14]), .IN2(n5), .IN3(data0[14]), .IN4(n4), .Q(
        data_o[14]) );
  AO22X1 U15 ( .IN1(data1[13]), .IN2(n5), .IN3(data0[13]), .IN4(n4), .Q(
        data_o[13]) );
  AO22X1 U16 ( .IN1(data1[12]), .IN2(n5), .IN3(data0[12]), .IN4(n4), .Q(
        data_o[12]) );
  AO22X1 U17 ( .IN1(data1[11]), .IN2(n5), .IN3(data0[11]), .IN4(n4), .Q(
        data_o[11]) );
  AO22X1 U18 ( .IN1(data1[10]), .IN2(n5), .IN3(data0[10]), .IN4(n4), .Q(
        data_o[10]) );
  AO22X1 U19 ( .IN1(data1[0]), .IN2(n5), .IN3(data0[0]), .IN4(n4), .Q(
        data_o[0]) );
  INVX0 U2 ( .INP(select1), .ZN(n1) );
  AND2X1 U3 ( .IN1(select0), .IN2(n1), .Q(n4) );
  NOR2X0 U20 ( .IN1(n1), .IN2(select0), .QN(n5) );
endmodule



    module node3_NODE_X0_NODE_Y3I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__ ( 
        \clk.clk , \reset.reset , \local_node.clk , 
        \local_node.buffer_full_in , \local_node.buffer_full_out , 
        \local_node.receiving_data , \local_node.sending_data , 
        \local_node.data_in , \local_node.data_out , \node_0.clk , 
        \node_0.buffer_full_in , \node_0.buffer_full_out , 
        \node_0.receiving_data , \node_0.sending_data , \node_0.data_in , 
        \node_0.data_out , \node_1.clk , \node_1.buffer_full_in , 
        \node_1.buffer_full_out , \node_1.receiving_data , 
        \node_1.sending_data , \node_1.data_in , \node_1.data_out  );
  input [15:0] \local_node.data_in ;
  output [15:0] \local_node.data_out ;
  input [15:0] \node_0.data_in ;
  output [15:0] \node_0.data_out ;
  input [15:0] \node_1.data_in ;
  output [15:0] \node_1.data_out ;
  input \clk.clk , \reset.reset , \local_node.buffer_full_in ,
         \local_node.receiving_data , \node_0.buffer_full_in ,
         \node_0.receiving_data , \node_1.buffer_full_in ,
         \node_1.receiving_data ;
  output \local_node.buffer_full_out , \local_node.sending_data ,
         \node_0.buffer_full_out , \node_0.sending_data ,
         \node_1.buffer_full_out , \node_1.sending_data ;
  inout \local_node.clk ,  \node_0.clk ,  \node_1.clk ;
  wire   \buffer_out[2][15] , \buffer_out[2][14] , \buffer_out[2][13] ,
         \buffer_out[2][12] , \buffer_out[2][11] , \buffer_out[2][10] ,
         \buffer_out[2][9] , \buffer_out[2][8] , \buffer_out[2][7] ,
         \buffer_out[2][6] , \buffer_out[2][5] , \buffer_out[2][4] ,
         \buffer_out[2][3] , \buffer_out[2][2] , \buffer_out[2][1] ,
         \buffer_out[2][0] , \buffer_out[1][15] , \buffer_out[1][14] ,
         \buffer_out[1][13] , \buffer_out[1][12] , \buffer_out[1][11] ,
         \buffer_out[1][10] , \buffer_out[1][9] , \buffer_out[1][8] ,
         \buffer_out[1][7] , \buffer_out[1][6] , \buffer_out[1][5] ,
         \buffer_out[1][4] , \buffer_out[1][3] , \buffer_out[1][2] ,
         \buffer_out[1][1] , \buffer_out[1][0] , \buffer_out[0][15] ,
         \buffer_out[0][14] , \buffer_out[0][13] , \buffer_out[0][12] ,
         \buffer_out[0][11] , \buffer_out[0][10] , \buffer_out[0][9] ,
         \buffer_out[0][8] , \buffer_out[0][7] , \buffer_out[0][6] ,
         \buffer_out[0][5] , \buffer_out[0][4] , \buffer_out[0][3] ,
         \buffer_out[0][2] , \buffer_out[0][1] , \buffer_out[0][0] ,
         \next_buffer_out[2][15] , \next_buffer_out[2][14] ,
         \next_buffer_out[2][13] , \next_buffer_out[2][12] ,
         \next_buffer_out[2][11] , \next_buffer_out[2][10] ,
         \next_buffer_out[2][9] , \next_buffer_out[2][8] ,
         \next_buffer_out[2][7] , \next_buffer_out[2][6] ,
         \next_buffer_out[2][5] , \next_buffer_out[2][4] ,
         \next_buffer_out[2][3] , \next_buffer_out[2][2] ,
         \next_buffer_out[2][1] , \next_buffer_out[2][0] ,
         \next_buffer_out[1][15] , \next_buffer_out[1][14] ,
         \next_buffer_out[1][13] , \next_buffer_out[1][12] ,
         \next_buffer_out[1][11] , \next_buffer_out[1][10] ,
         \next_buffer_out[1][9] , \next_buffer_out[1][8] ,
         \next_buffer_out[1][7] , \next_buffer_out[1][6] ,
         \next_buffer_out[1][5] , \next_buffer_out[1][4] ,
         \next_buffer_out[1][3] , \next_buffer_out[1][2] ,
         \next_buffer_out[1][1] , \next_buffer_out[1][0] ,
         \next_buffer_out[0][15] , \next_buffer_out[0][14] ,
         \next_buffer_out[0][13] , \next_buffer_out[0][12] ,
         \next_buffer_out[0][11] , \next_buffer_out[0][10] ,
         \next_buffer_out[0][9] , \next_buffer_out[0][8] ,
         \next_buffer_out[0][7] , \next_buffer_out[0][6] ,
         \next_buffer_out[0][5] , \next_buffer_out[0][4] ,
         \next_buffer_out[0][3] , \next_buffer_out[0][2] ,
         \next_buffer_out[0][1] , \next_buffer_out[0][0] ;
  wire   [2:0] buffer_full_in;
  wire   [2:0] receiving_data;
  wire   [2:0] pop_v;
  wire   [2:0] data_valid;
  wire   [2:0] next_data_valid;
  wire   [1:0] grant_1;
  wire   [1:0] grant_2;
  tri   \local_node.buffer_full_in ;
  tri   \local_node.buffer_full_out ;
  tri   \local_node.receiving_data ;
  tri   \local_node.sending_data ;
  tri   [15:0] \local_node.data_in ;
  tri   [15:0] \local_node.data_out ;

  converter_out_I_n_node_interface_dut_ c2 ( .\n.buffer_full_in (
        \local_node.buffer_full_in ), .\n.receiving_data (
        \local_node.receiving_data ), .\n.data_in (\local_node.data_in ), 
        .\n.buffer_full_out (\local_node.buffer_full_out ), .\n.sending_data (
        \local_node.sending_data ), .\n.data_out (\local_node.data_out ), 
        .buffer_full_in(1'b0), .receiving_data(1'b0), .data_in({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  fifo_kev_57 \genblk1[0].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[0]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[0]), .data_out({\buffer_out[0][15] , 
        \buffer_out[0][14] , \buffer_out[0][13] , \buffer_out[0][12] , 
        \buffer_out[0][11] , \buffer_out[0][10] , \buffer_out[0][9] , 
        \buffer_out[0][8] , \buffer_out[0][7] , \buffer_out[0][6] , 
        \buffer_out[0][5] , \buffer_out[0][4] , \buffer_out[0][3] , 
        \buffer_out[0][2] , \buffer_out[0][1] , \buffer_out[0][0] }), 
        .next_data_out({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] , 
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .next_data_valid(
        next_data_valid[0]) );
  address_counter_57 \genblk1[0].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] }), 
        .buffer_data_valid(next_data_valid[0]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .buffer_pop(
        pop_v[0]), .receiving_data(1'b0) );
  fifo_kev_56 \genblk1[1].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[1]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[1]), .data_out({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), 
        .next_data_out({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] , 
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .next_data_valid(
        next_data_valid[1]) );
  address_counter_56 \genblk1[1].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] }), 
        .buffer_data_valid(next_data_valid[1]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .buffer_pop(
        pop_v[1]), .receiving_data(1'b0) );
  fifo_kev_55 \genblk1[2].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[2]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[2]), .data_out({\buffer_out[2][15] , 
        \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] , 
        \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] , 
        \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] , 
        \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] , 
        \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] }), 
        .next_data_out({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] , 
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .next_data_valid(
        next_data_valid[2]) );
  address_counter_55 \genblk1[2].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] }), 
        .buffer_data_valid(next_data_valid[2]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .buffer_pop(
        pop_v[2]), .receiving_data(1'b0) );
  converter_in_I_n_node_interface_dut__22 \genblk2.c0  ( .\n.buffer_full_in (
        \node_0.buffer_full_in ), .\n.receiving_data (\node_0.receiving_data ), 
        .\n.data_in (\node_0.data_in ), .\n.buffer_full_out (
        \node_0.buffer_full_out ), .\n.sending_data (\node_0.sending_data ), 
        .\n.data_out (\node_0.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_in_I_n_node_interface_dut__21 \genblk2.c1  ( .\n.buffer_full_in (
        \node_1.buffer_full_in ), .\n.receiving_data (\node_1.receiving_data ), 
        .\n.data_in (\node_1.data_in ), .\n.buffer_full_out (
        \node_1.buffer_full_out ), .\n.sending_data (\node_1.sending_data ), 
        .\n.data_out (\node_1.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  controller3_sw \genblk2.sw  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .packet_addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .local_addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b1, 1'b1}), .packet_valid(data_valid), .buffer_full_in({1'b0, 1'b0, 
        1'b0}), .grant_1(grant_1), .grant_2(grant_2), .pop_v(pop_v) );
  mux2_1_19 \genblk2.mux_e  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[2][15] , 
        \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] , 
        \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] , 
        \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] , 
        \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] , 
        \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] }), 
        .select0(grant_1[0]), .select1(grant_1[1]) );
  mux2_1_18 \genblk2.mux_l  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), 
        .select0(grant_2[0]), .select1(grant_2[1]) );
endmodule


module fifo_kev_54 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_109 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_54 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_109 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_108 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_54 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_108 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_54_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_54 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_54 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_54 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_54_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_53 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_107 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_53 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_107 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_106 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_53 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_106 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_53_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_53 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_53 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_53 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_53_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_52 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_105 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_52 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_105 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_104 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_52 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_104 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_52_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_52 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_52 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_52 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_52_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module converter_in_I_n_node_interface_dut__20 ( \n.buffer_full_in , 
        \n.receiving_data , \n.data_in , \n.buffer_full_out , \n.sending_data , 
        \n.data_out , buffer_full_out, sending_data, data_out, buffer_full_in, 
        receiving_data, data_in );
  input [15:0] \n.data_in ;
  output [15:0] \n.data_out ;
  output [15:0] data_out;
  input [15:0] data_in;
  input \n.buffer_full_in , \n.receiving_data , buffer_full_in, receiving_data;
  output \n.buffer_full_out , \n.sending_data , buffer_full_out, sending_data;
  wire   \n.buffer_full_in , \n.receiving_data , buffer_full_in,
         receiving_data;
  assign buffer_full_out = \n.buffer_full_in ;
  assign sending_data = \n.receiving_data ;
  assign data_out[15] = \n.data_in  [15];
  assign data_out[14] = \n.data_in  [14];
  assign data_out[13] = \n.data_in  [13];
  assign data_out[12] = \n.data_in  [12];
  assign data_out[11] = \n.data_in  [11];
  assign data_out[10] = \n.data_in  [10];
  assign data_out[9] = \n.data_in  [9];
  assign data_out[8] = \n.data_in  [8];
  assign data_out[7] = \n.data_in  [7];
  assign data_out[6] = \n.data_in  [6];
  assign data_out[5] = \n.data_in  [5];
  assign data_out[4] = \n.data_in  [4];
  assign data_out[3] = \n.data_in  [3];
  assign data_out[2] = \n.data_in  [2];
  assign data_out[1] = \n.data_in  [1];
  assign data_out[0] = \n.data_in  [0];
  assign \n.buffer_full_out  = buffer_full_in;
  assign \n.sending_data  = receiving_data;
  assign \n.data_out  [15] = data_in[15];
  assign \n.data_out  [14] = data_in[14];
  assign \n.data_out  [13] = data_in[13];
  assign \n.data_out  [12] = data_in[12];
  assign \n.data_out  [11] = data_in[11];
  assign \n.data_out  [10] = data_in[10];
  assign \n.data_out  [9] = data_in[9];
  assign \n.data_out  [8] = data_in[8];
  assign \n.data_out  [7] = data_in[7];
  assign \n.data_out  [6] = data_in[6];
  assign \n.data_out  [5] = data_in[5];
  assign \n.data_out  [4] = data_in[4];
  assign \n.data_out  [3] = data_in[3];
  assign \n.data_out  [2] = data_in[2];
  assign \n.data_out  [1] = data_in[1];
  assign \n.data_out  [0] = data_in[0];

endmodule


module flipflop_BITS2_17 ( clk, data_i, data_o );
  input [1:0] data_i;
  output [1:0] data_o;
  input clk;


  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS2_17 ( clk, enable_i, reset, data_i, data_o );
  input [1:0] data_i;
  input [1:0] data_o;
  input clk, enable_i, reset;
  wire   n10, n11, n1, n5, n7, n8, n9;
  wire   [1:0] write_data;

  AOI22X1 U5 ( .IN1(enable_i), .IN2(data_i[1]), .IN3(n10), .IN4(n1), .QN(n9)
         );
  AOI22X1 U6 ( .IN1(data_i[0]), .IN2(enable_i), .IN3(n11), .IN4(n1), .QN(n8)
         );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n9), .QN(write_data[1]) );
  NOR2X0 U4 ( .IN1(reset), .IN2(n8), .QN(write_data[0]) );
  AND2X1 U7 ( .IN1(data_o[1]), .IN2(n7), .Q(n10) );
  AND2X1 U8 ( .IN1(data_o[0]), .IN2(n5), .Q(n11) );
  flipflop_BITS2_17 FF ( .clk(clk), .data_i(write_data), .data_o({n7, n5}) );
endmodule


module flipflop_BITS1_81 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_81 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_81 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter2_17 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [1:0] request;
  output [1:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   tail_en, n1, n2;
  wire   [1:0] req_i;
  wire   [1:0] req_o;

  AND3X1 U10 ( .IN1(request[1]), .IN2(n1), .IN3(n2), .Q(grant[1]) );
  AND3X1 U11 ( .IN1(request[0]), .IN2(n2), .IN3(request[1]), .Q(tail_en) );
  INVX0 U6 ( .INP(request[0]), .ZN(n1) );
  NOR2X0 U7 ( .IN1(buffer_full_i), .IN2(n1), .QN(grant[0]) );
  INVX0 U8 ( .INP(buffer_full_i), .ZN(n2) );
  OA21X1 U9 ( .IN1(request[1]), .IN2(request[0]), .IN3(n2), .Q(grant_v_o) );
  register_BITS2_17 req_record ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i({1'b1, 1'b0}), .data_o({1'b0, 1'b0}) );
  register_BITS1_81 tail ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i(1'b1), .data_o(1'b0) );
endmodule


module flipflop_BITS2_16 ( clk, data_i, data_o );
  input [1:0] data_i;
  output [1:0] data_o;
  input clk;


  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS2_16 ( clk, enable_i, reset, data_i, data_o );
  input [1:0] data_i;
  input [1:0] data_o;
  input clk, enable_i, reset;
  wire   n10, n11, n1, n5, n7, n8, n9;
  wire   [1:0] write_data;

  AOI22X1 U5 ( .IN1(enable_i), .IN2(data_i[1]), .IN3(n10), .IN4(n1), .QN(n9)
         );
  AOI22X1 U6 ( .IN1(data_i[0]), .IN2(enable_i), .IN3(n11), .IN4(n1), .QN(n8)
         );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n9), .QN(write_data[1]) );
  NOR2X0 U4 ( .IN1(reset), .IN2(n8), .QN(write_data[0]) );
  AND2X1 U7 ( .IN1(data_o[1]), .IN2(n7), .Q(n10) );
  AND2X1 U8 ( .IN1(data_o[0]), .IN2(n5), .Q(n11) );
  flipflop_BITS2_16 FF ( .clk(clk), .data_i(write_data), .data_o({n7, n5}) );
endmodule


module flipflop_BITS1_80 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_80 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_80 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter2_16 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [1:0] request;
  output [1:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   tail_en, n1, n2;
  wire   [1:0] req_i;
  wire   [1:0] req_o;

  AND3X1 U10 ( .IN1(request[1]), .IN2(n1), .IN3(n2), .Q(grant[1]) );
  AND3X1 U11 ( .IN1(request[0]), .IN2(n2), .IN3(request[1]), .Q(tail_en) );
  INVX0 U6 ( .INP(request[0]), .ZN(n1) );
  NOR2X0 U7 ( .IN1(buffer_full_i), .IN2(n1), .QN(grant[0]) );
  INVX0 U8 ( .INP(buffer_full_i), .ZN(n2) );
  OA21X1 U9 ( .IN1(request[1]), .IN2(request[0]), .IN3(n2), .Q(grant_v_o) );
  register_BITS2_16 req_record ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i({1'b1, 1'b0}), .data_o({1'b0, 1'b0}) );
  register_BITS1_80 tail ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i(1'b1), .data_o(1'b0) );
endmodule


module dccl_54 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_53 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_52 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module controller3_se ( clk, rst, .packet_addr({\packet_addr[2][7] , 
        \packet_addr[2][6] , \packet_addr[2][5] , \packet_addr[2][4] , 
        \packet_addr[2][3] , \packet_addr[2][2] , \packet_addr[2][1] , 
        \packet_addr[2][0] , \packet_addr[1][7] , \packet_addr[1][6] , 
        \packet_addr[1][5] , \packet_addr[1][4] , \packet_addr[1][3] , 
        \packet_addr[1][2] , \packet_addr[1][1] , \packet_addr[1][0] , 
        \packet_addr[0][7] , \packet_addr[0][6] , \packet_addr[0][5] , 
        \packet_addr[0][4] , \packet_addr[0][3] , \packet_addr[0][2] , 
        \packet_addr[0][1] , \packet_addr[0][0] }), local_addr, packet_valid, 
        buffer_full_in, grant_1, grant_2, grant_v, pop_v );
  input [7:0] local_addr;
  input [2:0] packet_valid;
  input [2:0] buffer_full_in;
  output [1:0] grant_1;
  output [1:0] grant_2;
  output [2:0] grant_v;
  output [2:0] pop_v;
  input clk, rst, \packet_addr[2][7] , \packet_addr[2][6] ,
         \packet_addr[2][5] , \packet_addr[2][4] , \packet_addr[2][3] ,
         \packet_addr[2][2] , \packet_addr[2][1] , \packet_addr[2][0] ,
         \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] ,
         \packet_addr[1][4] , \packet_addr[1][3] , \packet_addr[1][2] ,
         \packet_addr[1][1] , \packet_addr[1][0] , \packet_addr[0][7] ,
         \packet_addr[0][6] , \packet_addr[0][5] , \packet_addr[0][4] ,
         \packet_addr[0][3] , \packet_addr[0][2] , \packet_addr[0][1] ,
         \packet_addr[0][0] ;
  wire   \grant_2[1] , \request[2][1] , \request[2][0] , \request[1][1] ,
         \request[1][0] , \request[0][0] , n1;
  assign pop_v[1] = \grant_2[1] ;
  assign grant_2[1] = \grant_2[1] ;

  OR2X1 U3 ( .IN1(grant_v[0]), .IN2(grant_1[1]), .Q(pop_v[2]) );
  OR2X1 U4 ( .IN1(grant_1[0]), .IN2(grant_2[0]), .Q(pop_v[0]) );
  NOR2X0 U1 ( .IN1(n1), .IN2(buffer_full_in[0]), .QN(grant_v[0]) );
  INVX0 U2 ( .INP(\request[0][0] ), .ZN(n1) );
  arbiter2_17 arbiter_w ( .clk(clk), .rst(rst), .request({\request[1][1] , 
        \request[1][0] }), .buffer_full_i(buffer_full_in[1]), .grant(grant_1), 
        .grant_v_o(grant_v[1]) );
  arbiter2_16 arbiter_l ( .clk(clk), .rst(rst), .request({\request[2][1] , 
        \request[2][0] }), .buffer_full_i(buffer_full_in[2]), .grant({
        \grant_2[1] , grant_2[0]}), .grant_v_o(grant_v[2]) );
  dccl_54 dccl_n ( .packet_addr_y_i({\packet_addr[0][3] , \packet_addr[0][2] , 
        \packet_addr[0][1] , \packet_addr[0][0] }), .packet_addr_x_i({
        \packet_addr[0][7] , \packet_addr[0][6] , \packet_addr[0][5] , 
        \packet_addr[0][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[0]), 
        .west_req(\request[1][0] ), .local_req(\request[2][0] ) );
  dccl_53 dccl_w ( .packet_addr_y_i({\packet_addr[1][3] , \packet_addr[1][2] , 
        \packet_addr[1][1] , \packet_addr[1][0] }), .packet_addr_x_i({
        \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] , 
        \packet_addr[1][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[1]), 
        .local_req(\request[2][1] ) );
  dccl_52 dccl_l ( .packet_addr_y_i({\packet_addr[2][3] , \packet_addr[2][2] , 
        \packet_addr[2][1] , \packet_addr[2][0] }), .packet_addr_x_i({
        \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] , 
        \packet_addr[2][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[2]), 
        .north_req(\request[0][0] ), .west_req(\request[1][1] ) );
endmodule


module mux2_1_17 ( data0, data1, select0, select1, data_o );
  input [15:0] data0;
  input [15:0] data1;
  output [15:0] data_o;
  input select0, select1;
  wire   n1, n4, n5;

  AO22X1 U4 ( .IN1(data1[9]), .IN2(n5), .IN3(data0[9]), .IN4(n4), .Q(data_o[9]) );
  AO22X1 U5 ( .IN1(data1[8]), .IN2(n5), .IN3(data0[8]), .IN4(n4), .Q(data_o[8]) );
  AO22X1 U6 ( .IN1(data1[7]), .IN2(n5), .IN3(data0[7]), .IN4(n4), .Q(data_o[7]) );
  AO22X1 U7 ( .IN1(data1[6]), .IN2(n5), .IN3(data0[6]), .IN4(n4), .Q(data_o[6]) );
  AO22X1 U8 ( .IN1(data1[5]), .IN2(n5), .IN3(data0[5]), .IN4(n4), .Q(data_o[5]) );
  AO22X1 U9 ( .IN1(data1[4]), .IN2(n5), .IN3(data0[4]), .IN4(n4), .Q(data_o[4]) );
  AO22X1 U10 ( .IN1(data1[3]), .IN2(n5), .IN3(data0[3]), .IN4(n4), .Q(
        data_o[3]) );
  AO22X1 U11 ( .IN1(data1[2]), .IN2(n5), .IN3(data0[2]), .IN4(n4), .Q(
        data_o[2]) );
  AO22X1 U12 ( .IN1(data1[1]), .IN2(n5), .IN3(data0[1]), .IN4(n4), .Q(
        data_o[1]) );
  AO22X1 U13 ( .IN1(data1[15]), .IN2(n5), .IN3(data0[15]), .IN4(n4), .Q(
        data_o[15]) );
  AO22X1 U14 ( .IN1(data1[14]), .IN2(n5), .IN3(data0[14]), .IN4(n4), .Q(
        data_o[14]) );
  AO22X1 U15 ( .IN1(data1[13]), .IN2(n5), .IN3(data0[13]), .IN4(n4), .Q(
        data_o[13]) );
  AO22X1 U16 ( .IN1(data1[12]), .IN2(n5), .IN3(data0[12]), .IN4(n4), .Q(
        data_o[12]) );
  AO22X1 U17 ( .IN1(data1[11]), .IN2(n5), .IN3(data0[11]), .IN4(n4), .Q(
        data_o[11]) );
  AO22X1 U18 ( .IN1(data1[10]), .IN2(n5), .IN3(data0[10]), .IN4(n4), .Q(
        data_o[10]) );
  AO22X1 U19 ( .IN1(data1[0]), .IN2(n5), .IN3(data0[0]), .IN4(n4), .Q(
        data_o[0]) );
  INVX0 U2 ( .INP(select1), .ZN(n1) );
  AND2X1 U3 ( .IN1(select0), .IN2(n1), .Q(n4) );
  NOR2X0 U20 ( .IN1(n1), .IN2(select0), .QN(n5) );
endmodule


module mux2_1_16 ( data0, data1, select0, select1, data_o );
  input [15:0] data0;
  input [15:0] data1;
  output [15:0] data_o;
  input select0, select1;
  wire   n1, n4, n5;

  AO22X1 U4 ( .IN1(data1[9]), .IN2(n5), .IN3(data0[9]), .IN4(n4), .Q(data_o[9]) );
  AO22X1 U5 ( .IN1(data1[8]), .IN2(n5), .IN3(data0[8]), .IN4(n4), .Q(data_o[8]) );
  AO22X1 U6 ( .IN1(data1[7]), .IN2(n5), .IN3(data0[7]), .IN4(n4), .Q(data_o[7]) );
  AO22X1 U7 ( .IN1(data1[6]), .IN2(n5), .IN3(data0[6]), .IN4(n4), .Q(data_o[6]) );
  AO22X1 U8 ( .IN1(data1[5]), .IN2(n5), .IN3(data0[5]), .IN4(n4), .Q(data_o[5]) );
  AO22X1 U9 ( .IN1(data1[4]), .IN2(n5), .IN3(data0[4]), .IN4(n4), .Q(data_o[4]) );
  AO22X1 U10 ( .IN1(data1[3]), .IN2(n5), .IN3(data0[3]), .IN4(n4), .Q(
        data_o[3]) );
  AO22X1 U11 ( .IN1(data1[2]), .IN2(n5), .IN3(data0[2]), .IN4(n4), .Q(
        data_o[2]) );
  AO22X1 U12 ( .IN1(data1[1]), .IN2(n5), .IN3(data0[1]), .IN4(n4), .Q(
        data_o[1]) );
  AO22X1 U13 ( .IN1(data1[15]), .IN2(n5), .IN3(data0[15]), .IN4(n4), .Q(
        data_o[15]) );
  AO22X1 U14 ( .IN1(data1[14]), .IN2(n5), .IN3(data0[14]), .IN4(n4), .Q(
        data_o[14]) );
  AO22X1 U15 ( .IN1(data1[13]), .IN2(n5), .IN3(data0[13]), .IN4(n4), .Q(
        data_o[13]) );
  AO22X1 U16 ( .IN1(data1[12]), .IN2(n5), .IN3(data0[12]), .IN4(n4), .Q(
        data_o[12]) );
  AO22X1 U17 ( .IN1(data1[11]), .IN2(n5), .IN3(data0[11]), .IN4(n4), .Q(
        data_o[11]) );
  AO22X1 U18 ( .IN1(data1[10]), .IN2(n5), .IN3(data0[10]), .IN4(n4), .Q(
        data_o[10]) );
  AO22X1 U19 ( .IN1(data1[0]), .IN2(n5), .IN3(data0[0]), .IN4(n4), .Q(
        data_o[0]) );
  INVX0 U2 ( .INP(select1), .ZN(n1) );
  AND2X1 U3 ( .IN1(select0), .IN2(n1), .Q(n4) );
  NOR2X0 U20 ( .IN1(n1), .IN2(select0), .QN(n5) );
endmodule



    module node3_NODE_X3_NODE_Y3I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__ ( 
        \clk.clk , \reset.reset , \local_node.clk , 
        \local_node.buffer_full_in , \local_node.buffer_full_out , 
        \local_node.receiving_data , \local_node.sending_data , 
        \local_node.data_in , \local_node.data_out , \node_0.clk , 
        \node_0.buffer_full_in , \node_0.buffer_full_out , 
        \node_0.receiving_data , \node_0.sending_data , \node_0.data_in , 
        \node_0.data_out , \node_1.clk , \node_1.buffer_full_in , 
        \node_1.buffer_full_out , \node_1.receiving_data , 
        \node_1.sending_data , \node_1.data_in , \node_1.data_out  );
  input [15:0] \local_node.data_in ;
  output [15:0] \local_node.data_out ;
  input [15:0] \node_0.data_in ;
  output [15:0] \node_0.data_out ;
  input [15:0] \node_1.data_in ;
  output [15:0] \node_1.data_out ;
  input \clk.clk , \reset.reset , \local_node.buffer_full_in ,
         \local_node.receiving_data , \node_0.buffer_full_in ,
         \node_0.receiving_data , \node_1.buffer_full_in ,
         \node_1.receiving_data ;
  output \local_node.buffer_full_out , \local_node.sending_data ,
         \node_0.buffer_full_out , \node_0.sending_data ,
         \node_1.buffer_full_out , \node_1.sending_data ;
  inout \local_node.clk ,  \node_0.clk ,  \node_1.clk ;
  wire   \buffer_out[2][15] , \buffer_out[2][14] , \buffer_out[2][13] ,
         \buffer_out[2][12] , \buffer_out[2][11] , \buffer_out[2][10] ,
         \buffer_out[2][9] , \buffer_out[2][8] , \buffer_out[2][7] ,
         \buffer_out[2][6] , \buffer_out[2][5] , \buffer_out[2][4] ,
         \buffer_out[2][3] , \buffer_out[2][2] , \buffer_out[2][1] ,
         \buffer_out[2][0] , \buffer_out[1][15] , \buffer_out[1][14] ,
         \buffer_out[1][13] , \buffer_out[1][12] , \buffer_out[1][11] ,
         \buffer_out[1][10] , \buffer_out[1][9] , \buffer_out[1][8] ,
         \buffer_out[1][7] , \buffer_out[1][6] , \buffer_out[1][5] ,
         \buffer_out[1][4] , \buffer_out[1][3] , \buffer_out[1][2] ,
         \buffer_out[1][1] , \buffer_out[1][0] , \buffer_out[0][15] ,
         \buffer_out[0][14] , \buffer_out[0][13] , \buffer_out[0][12] ,
         \buffer_out[0][11] , \buffer_out[0][10] , \buffer_out[0][9] ,
         \buffer_out[0][8] , \buffer_out[0][7] , \buffer_out[0][6] ,
         \buffer_out[0][5] , \buffer_out[0][4] , \buffer_out[0][3] ,
         \buffer_out[0][2] , \buffer_out[0][1] , \buffer_out[0][0] ,
         \next_buffer_out[2][15] , \next_buffer_out[2][14] ,
         \next_buffer_out[2][13] , \next_buffer_out[2][12] ,
         \next_buffer_out[2][11] , \next_buffer_out[2][10] ,
         \next_buffer_out[2][9] , \next_buffer_out[2][8] ,
         \next_buffer_out[2][7] , \next_buffer_out[2][6] ,
         \next_buffer_out[2][5] , \next_buffer_out[2][4] ,
         \next_buffer_out[2][3] , \next_buffer_out[2][2] ,
         \next_buffer_out[2][1] , \next_buffer_out[2][0] ,
         \next_buffer_out[1][15] , \next_buffer_out[1][14] ,
         \next_buffer_out[1][13] , \next_buffer_out[1][12] ,
         \next_buffer_out[1][11] , \next_buffer_out[1][10] ,
         \next_buffer_out[1][9] , \next_buffer_out[1][8] ,
         \next_buffer_out[1][7] , \next_buffer_out[1][6] ,
         \next_buffer_out[1][5] , \next_buffer_out[1][4] ,
         \next_buffer_out[1][3] , \next_buffer_out[1][2] ,
         \next_buffer_out[1][1] , \next_buffer_out[1][0] ,
         \next_buffer_out[0][15] , \next_buffer_out[0][14] ,
         \next_buffer_out[0][13] , \next_buffer_out[0][12] ,
         \next_buffer_out[0][11] , \next_buffer_out[0][10] ,
         \next_buffer_out[0][9] , \next_buffer_out[0][8] ,
         \next_buffer_out[0][7] , \next_buffer_out[0][6] ,
         \next_buffer_out[0][5] , \next_buffer_out[0][4] ,
         \next_buffer_out[0][3] , \next_buffer_out[0][2] ,
         \next_buffer_out[0][1] , \next_buffer_out[0][0] ;
  wire   [2:0] buffer_full_in;
  wire   [2:0] receiving_data;
  wire   [2:0] pop_v;
  wire   [2:0] data_valid;
  wire   [2:0] next_data_valid;
  wire   [1:0] grant_1;
  wire   [1:0] grant_2;
  tri   \local_node.buffer_full_in ;
  tri   \local_node.buffer_full_out ;
  tri   \local_node.receiving_data ;
  tri   \local_node.sending_data ;
  tri   [15:0] \local_node.data_in ;
  tri   [15:0] \local_node.data_out ;

  converter_out_I_n_node_interface_dut_ c2 ( .\n.buffer_full_in (
        \local_node.buffer_full_in ), .\n.receiving_data (
        \local_node.receiving_data ), .\n.data_in (\local_node.data_in ), 
        .\n.buffer_full_out (\local_node.buffer_full_out ), .\n.sending_data (
        \local_node.sending_data ), .\n.data_out (\local_node.data_out ), 
        .buffer_full_in(1'b0), .receiving_data(1'b0), .data_in({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  fifo_kev_54 \genblk1[0].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[0]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[0]), .data_out({\buffer_out[0][15] , 
        \buffer_out[0][14] , \buffer_out[0][13] , \buffer_out[0][12] , 
        \buffer_out[0][11] , \buffer_out[0][10] , \buffer_out[0][9] , 
        \buffer_out[0][8] , \buffer_out[0][7] , \buffer_out[0][6] , 
        \buffer_out[0][5] , \buffer_out[0][4] , \buffer_out[0][3] , 
        \buffer_out[0][2] , \buffer_out[0][1] , \buffer_out[0][0] }), 
        .next_data_out({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] , 
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .next_data_valid(
        next_data_valid[0]) );
  address_counter_54 \genblk1[0].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] }), 
        .buffer_data_valid(next_data_valid[0]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .buffer_pop(
        pop_v[0]), .receiving_data(1'b0) );
  fifo_kev_53 \genblk1[1].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[1]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[1]), .data_out({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), 
        .next_data_out({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] , 
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .next_data_valid(
        next_data_valid[1]) );
  address_counter_53 \genblk1[1].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] }), 
        .buffer_data_valid(next_data_valid[1]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .buffer_pop(
        pop_v[1]), .receiving_data(1'b0) );
  fifo_kev_52 \genblk1[2].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[2]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[2]), .data_out({\buffer_out[2][15] , 
        \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] , 
        \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] , 
        \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] , 
        \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] , 
        \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] }), 
        .next_data_out({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] , 
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .next_data_valid(
        next_data_valid[2]) );
  address_counter_52 \genblk1[2].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] }), 
        .buffer_data_valid(next_data_valid[2]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .buffer_pop(
        pop_v[2]), .receiving_data(1'b0) );
  converter_in_I_n_node_interface_dut__20 \genblk2.c0  ( .\n.buffer_full_in (
        \node_0.buffer_full_in ), .\n.receiving_data (\node_0.receiving_data ), 
        .\n.data_in (\node_0.data_in ), .\n.buffer_full_out (
        \node_0.buffer_full_out ), .\n.sending_data (\node_0.sending_data ), 
        .\n.data_out (\node_0.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_out_I_n_node_interface_dut_ \genblk2.c1  ( .\n.buffer_full_in (
        \node_1.buffer_full_in ), .\n.receiving_data (\node_1.receiving_data ), 
        .\n.data_in (\node_1.data_in ), .\n.buffer_full_out (
        \node_1.buffer_full_out ), .\n.sending_data (\node_1.sending_data ), 
        .\n.data_out (\node_1.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  controller3_se \genblk2.se  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .packet_addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .local_addr({1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 
        1'b1, 1'b1}), .packet_valid(data_valid), .buffer_full_in({1'b0, 1'b0, 
        1'b0}), .grant_1(grant_1), .grant_2(grant_2), .pop_v(pop_v) );
  mux2_1_17 \genblk2.mux_w  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[2][15] , 
        \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] , 
        \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] , 
        \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] , 
        \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] , 
        \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] }), 
        .select0(grant_1[0]), .select1(grant_1[1]) );
  mux2_1_16 \genblk2.mux_l  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), 
        .select0(grant_2[0]), .select1(grant_2[1]) );
endmodule


module fifo_kev_51 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_103 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_51 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_103 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_102 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_51 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_102 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_51_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_51 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_51 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_51 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_51_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_50 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_101 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_50 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_101 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_100 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_50 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_100 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_50_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_50 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_50 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_50 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_50_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_49 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_99 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_49 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_99 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_98 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_49 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_98 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_49_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_49 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_49 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_49 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_49_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_48 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_97 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_48 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_97 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_96 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_48 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_96 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_48_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_48 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_48 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_48 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_48_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module converter_in_I_n_node_interface_dut__19 ( \n.buffer_full_in , 
        \n.receiving_data , \n.data_in , \n.buffer_full_out , \n.sending_data , 
        \n.data_out , buffer_full_out, sending_data, data_out, buffer_full_in, 
        receiving_data, data_in );
  input [15:0] \n.data_in ;
  output [15:0] \n.data_out ;
  output [15:0] data_out;
  input [15:0] data_in;
  input \n.buffer_full_in , \n.receiving_data , buffer_full_in, receiving_data;
  output \n.buffer_full_out , \n.sending_data , buffer_full_out, sending_data;
  wire   \n.buffer_full_in , \n.receiving_data , buffer_full_in,
         receiving_data;
  assign buffer_full_out = \n.buffer_full_in ;
  assign sending_data = \n.receiving_data ;
  assign data_out[15] = \n.data_in  [15];
  assign data_out[14] = \n.data_in  [14];
  assign data_out[13] = \n.data_in  [13];
  assign data_out[12] = \n.data_in  [12];
  assign data_out[11] = \n.data_in  [11];
  assign data_out[10] = \n.data_in  [10];
  assign data_out[9] = \n.data_in  [9];
  assign data_out[8] = \n.data_in  [8];
  assign data_out[7] = \n.data_in  [7];
  assign data_out[6] = \n.data_in  [6];
  assign data_out[5] = \n.data_in  [5];
  assign data_out[4] = \n.data_in  [4];
  assign data_out[3] = \n.data_in  [3];
  assign data_out[2] = \n.data_in  [2];
  assign data_out[1] = \n.data_in  [1];
  assign data_out[0] = \n.data_in  [0];
  assign \n.buffer_full_out  = buffer_full_in;
  assign \n.sending_data  = receiving_data;
  assign \n.data_out  [15] = data_in[15];
  assign \n.data_out  [14] = data_in[14];
  assign \n.data_out  [13] = data_in[13];
  assign \n.data_out  [12] = data_in[12];
  assign \n.data_out  [11] = data_in[11];
  assign \n.data_out  [10] = data_in[10];
  assign \n.data_out  [9] = data_in[9];
  assign \n.data_out  [8] = data_in[8];
  assign \n.data_out  [7] = data_in[7];
  assign \n.data_out  [6] = data_in[6];
  assign \n.data_out  [5] = data_in[5];
  assign \n.data_out  [4] = data_in[4];
  assign \n.data_out  [3] = data_in[3];
  assign \n.data_out  [2] = data_in[2];
  assign \n.data_out  [1] = data_in[1];
  assign \n.data_out  [0] = data_in[0];

endmodule


module flipflop_BITS3_39 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_39 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n10, n11, n12, n2, n3, n1, n5, n7, n9;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n2), .IN3(n10), .IN4(n3), .Q(write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n2), .IN3(n11), .IN4(n3), .Q(write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n2), .IN3(n12), .IN4(n3), .Q(write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n3) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n2) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n10) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n11) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n12) );
  flipflop_BITS3_39 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS3_38 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_38 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_38 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS1_79 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_79 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_79 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_78 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_78 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_78 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter3_19 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [2:0] request;
  output [2:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[1][2] , \req_i[1][1] , \req_i[1][0] , \req_i[0][2] ,
         \req_i[0][1] , tail_en, N99, N100, N101, N110, N111, N118, N119, N120,
         N121, n26, n27, n28, n29, n1, n2, n3, n4;
  wire   [1:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N99 = request[0];
  assign N100 = request[1];
  assign N101 = request[2];

  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(N111), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(N110), .Q(\req_i[0][1] ) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N121), .D(tail_en), .Q(req_en[0]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N120), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N119), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N118), .Q(grant[0]) );
  AND2X1 U20 ( .IN1(n26), .IN2(N101), .Q(n27) );
  OR3X1 U21 ( .IN1(n3), .IN2(N111), .IN3(n28), .Q(N121) );
  NOR3X0 U22 ( .IN1(N99), .IN2(N100), .IN3(n28), .QN(N120) );
  NOR3X0 U23 ( .IN1(n2), .IN2(N99), .IN3(n28), .QN(N119) );
  NAND3X0 U24 ( .IN1(n2), .IN2(n3), .IN3(n1), .QN(n29) );
  AO22X1 U25 ( .IN1(N100), .IN2(N101), .IN3(N99), .IN4(N101), .Q(N111) );
  INVX0 U10 ( .INP(N101), .ZN(n3) );
  NAND2X1 U11 ( .IN1(n29), .IN2(n4), .QN(n28) );
  INVX0 U12 ( .INP(N99), .ZN(n1) );
  INVX0 U13 ( .INP(N100), .ZN(n2) );
  INVX0 U14 ( .INP(buffer_full_i), .ZN(n4) );
  NAND2X1 U15 ( .IN1(n1), .IN2(n2), .QN(n26) );
  NOR2X0 U16 ( .IN1(n1), .IN2(n28), .QN(N118) );
  NOR2X0 U17 ( .IN1(n1), .IN2(n2), .QN(N110) );
  OA21X1 U18 ( .IN1(N110), .IN2(n27), .IN3(n4), .Q(tail_en) );
  OA21X1 U19 ( .IN1(N101), .IN2(n26), .IN3(n4), .Q(grant_v_o) );
  register_BITS3_39 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][2] , \req_i[0][1] , 1'b0}), .data_o({
        1'b0, 1'b0, 1'b0}) );
  register_BITS3_38 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][2] , \req_i[1][1] , \req_i[1][0] }), 
        .data_o({1'b0, 1'b0, 1'b0}) );
  register_BITS1_79 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b1), .data_o(1'b0) );
  register_BITS1_78 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module flipflop_BITS3_37 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_37 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_37 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS3_36 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_36 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_36 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS1_77 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_77 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_77 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_76 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_76 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_76 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter3_18 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [2:0] request;
  output [2:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[1][2] , \req_i[1][1] , \req_i[1][0] , \req_i[0][2] ,
         \req_i[0][1] , tail_en, N99, N100, N101, N110, N111, N118, N119, N120,
         N121, n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [1:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N99 = request[0];
  assign N100 = request[1];
  assign N101 = request[2];

  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(N111), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(N110), .Q(\req_i[0][1] ) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N121), .D(tail_en), .Q(req_en[0]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N120), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N119), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N118), .Q(grant[0]) );
  AND2X1 U20 ( .IN1(n8), .IN2(N101), .Q(n7) );
  OR3X1 U21 ( .IN1(n3), .IN2(N111), .IN3(n6), .Q(N121) );
  NOR3X0 U22 ( .IN1(N99), .IN2(N100), .IN3(n6), .QN(N120) );
  NOR3X0 U23 ( .IN1(n2), .IN2(N99), .IN3(n6), .QN(N119) );
  NAND3X0 U24 ( .IN1(n2), .IN2(n3), .IN3(n1), .QN(n5) );
  AO22X1 U25 ( .IN1(N100), .IN2(N101), .IN3(N99), .IN4(N101), .Q(N111) );
  INVX0 U10 ( .INP(N101), .ZN(n3) );
  NAND2X1 U11 ( .IN1(n5), .IN2(n4), .QN(n6) );
  INVX0 U12 ( .INP(N99), .ZN(n1) );
  INVX0 U13 ( .INP(N100), .ZN(n2) );
  INVX0 U14 ( .INP(buffer_full_i), .ZN(n4) );
  NAND2X1 U15 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NOR2X0 U16 ( .IN1(n1), .IN2(n6), .QN(N118) );
  NOR2X0 U17 ( .IN1(n1), .IN2(n2), .QN(N110) );
  OA21X1 U18 ( .IN1(N110), .IN2(n7), .IN3(n4), .Q(tail_en) );
  OA21X1 U19 ( .IN1(N101), .IN2(n8), .IN3(n4), .Q(grant_v_o) );
  register_BITS3_37 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][2] , \req_i[0][1] , 1'b0}), .data_o({
        1'b0, 1'b0, 1'b0}) );
  register_BITS3_36 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][2] , \req_i[1][1] , \req_i[1][0] }), 
        .data_o({1'b0, 1'b0, 1'b0}) );
  register_BITS1_77 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b1), .data_o(1'b0) );
  register_BITS1_76 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module flipflop_BITS3_35 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_35 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_35 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS3_34 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_34 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_34 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS1_75 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_75 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_75 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_74 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_74 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_74 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter3_17 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [2:0] request;
  output [2:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[1][2] , \req_i[1][1] , \req_i[1][0] , \req_i[0][2] ,
         \req_i[0][1] , tail_en, N99, N100, N101, N110, N111, N118, N119, N120,
         N121, n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [1:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N99 = request[0];
  assign N100 = request[1];
  assign N101 = request[2];

  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(N111), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(N110), .Q(\req_i[0][1] ) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N121), .D(tail_en), .Q(req_en[0]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N120), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N119), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N118), .Q(grant[0]) );
  AND2X1 U20 ( .IN1(n8), .IN2(N101), .Q(n7) );
  OR3X1 U21 ( .IN1(n3), .IN2(N111), .IN3(n6), .Q(N121) );
  NOR3X0 U22 ( .IN1(N99), .IN2(N100), .IN3(n6), .QN(N120) );
  NOR3X0 U23 ( .IN1(n2), .IN2(N99), .IN3(n6), .QN(N119) );
  NAND3X0 U24 ( .IN1(n2), .IN2(n3), .IN3(n1), .QN(n5) );
  AO22X1 U25 ( .IN1(N100), .IN2(N101), .IN3(N99), .IN4(N101), .Q(N111) );
  INVX0 U10 ( .INP(N101), .ZN(n3) );
  NAND2X1 U11 ( .IN1(n5), .IN2(n4), .QN(n6) );
  INVX0 U12 ( .INP(N99), .ZN(n1) );
  INVX0 U13 ( .INP(N100), .ZN(n2) );
  INVX0 U14 ( .INP(buffer_full_i), .ZN(n4) );
  NAND2X1 U15 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NOR2X0 U16 ( .IN1(n1), .IN2(n6), .QN(N118) );
  NOR2X0 U17 ( .IN1(n1), .IN2(n2), .QN(N110) );
  OA21X1 U18 ( .IN1(N110), .IN2(n7), .IN3(n4), .Q(tail_en) );
  OA21X1 U19 ( .IN1(N101), .IN2(n8), .IN3(n4), .Q(grant_v_o) );
  register_BITS3_35 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][2] , \req_i[0][1] , 1'b0}), .data_o({
        1'b0, 1'b0, 1'b0}) );
  register_BITS3_34 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][2] , \req_i[1][1] , \req_i[1][0] }), 
        .data_o({1'b0, 1'b0, 1'b0}) );
  register_BITS1_75 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b1), .data_o(1'b0) );
  register_BITS1_74 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module dccl_51 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_50 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_49 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_48 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module controller4_edge_n_1 ( clk, rst, .packet_addr({\packet_addr[3][7] , 
        \packet_addr[3][6] , \packet_addr[3][5] , \packet_addr[3][4] , 
        \packet_addr[3][3] , \packet_addr[3][2] , \packet_addr[3][1] , 
        \packet_addr[3][0] , \packet_addr[2][7] , \packet_addr[2][6] , 
        \packet_addr[2][5] , \packet_addr[2][4] , \packet_addr[2][3] , 
        \packet_addr[2][2] , \packet_addr[2][1] , \packet_addr[2][0] , 
        \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] , 
        \packet_addr[1][4] , \packet_addr[1][3] , \packet_addr[1][2] , 
        \packet_addr[1][1] , \packet_addr[1][0] , \packet_addr[0][7] , 
        \packet_addr[0][6] , \packet_addr[0][5] , \packet_addr[0][4] , 
        \packet_addr[0][3] , \packet_addr[0][2] , \packet_addr[0][1] , 
        \packet_addr[0][0] }), local_addr, packet_valid, buffer_full_in, 
        grant_1, grant_2, grant_3, grant_v, pop_v );
  input [7:0] local_addr;
  input [3:0] packet_valid;
  input [3:0] buffer_full_in;
  output [2:0] grant_1;
  output [2:0] grant_2;
  output [2:0] grant_3;
  output [3:0] grant_v;
  output [3:0] pop_v;
  input clk, rst, \packet_addr[3][7] , \packet_addr[3][6] ,
         \packet_addr[3][5] , \packet_addr[3][4] , \packet_addr[3][3] ,
         \packet_addr[3][2] , \packet_addr[3][1] , \packet_addr[3][0] ,
         \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] ,
         \packet_addr[2][4] , \packet_addr[2][3] , \packet_addr[2][2] ,
         \packet_addr[2][1] , \packet_addr[2][0] , \packet_addr[1][7] ,
         \packet_addr[1][6] , \packet_addr[1][5] , \packet_addr[1][4] ,
         \packet_addr[1][3] , \packet_addr[1][2] , \packet_addr[1][1] ,
         \packet_addr[1][0] , \packet_addr[0][7] , \packet_addr[0][6] ,
         \packet_addr[0][5] , \packet_addr[0][4] , \packet_addr[0][3] ,
         \packet_addr[0][2] , \packet_addr[0][1] , \packet_addr[0][0] ;
  wire   \request[3][2] , \request[3][1] , \request[3][0] , \request[2][2] ,
         \request[2][1] , \request[2][0] , \request[1][2] , \request[1][1] ,
         \request[1][0] , \request[0][0] , n1;

  OR3X1 U3 ( .IN1(grant_2[2]), .IN2(grant_1[2]), .IN3(grant_v[0]), .Q(pop_v[3]) );
  OR2X1 U4 ( .IN1(grant_1[1]), .IN2(grant_3[2]), .Q(pop_v[2]) );
  OR2X1 U5 ( .IN1(grant_2[1]), .IN2(grant_3[1]), .Q(pop_v[1]) );
  OR3X1 U6 ( .IN1(grant_3[0]), .IN2(grant_2[0]), .IN3(grant_1[0]), .Q(pop_v[0]) );
  NOR2X0 U1 ( .IN1(n1), .IN2(buffer_full_in[0]), .QN(grant_v[0]) );
  INVX0 U2 ( .INP(\request[0][0] ), .ZN(n1) );
  arbiter3_19 arbiter_e ( .clk(clk), .rst(rst), .request({\request[1][2] , 
        \request[1][1] , \request[1][0] }), .buffer_full_i(buffer_full_in[1]), 
        .grant(grant_1), .grant_v_o(grant_v[1]) );
  arbiter3_18 arbiter_w ( .clk(clk), .rst(rst), .request({\request[2][2] , 
        \request[2][1] , \request[2][0] }), .buffer_full_i(buffer_full_in[2]), 
        .grant(grant_2), .grant_v_o(grant_v[2]) );
  arbiter3_17 arbiter_l ( .clk(clk), .rst(rst), .request({\request[3][2] , 
        \request[3][1] , \request[3][0] }), .buffer_full_i(buffer_full_in[3]), 
        .grant(grant_3), .grant_v_o(grant_v[3]) );
  dccl_51 dccl_s ( .packet_addr_y_i({\packet_addr[0][3] , \packet_addr[0][2] , 
        \packet_addr[0][1] , \packet_addr[0][0] }), .packet_addr_x_i({
        \packet_addr[0][7] , \packet_addr[0][6] , \packet_addr[0][5] , 
        \packet_addr[0][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[0]), 
        .east_req(\request[1][0] ), .west_req(\request[2][0] ), .local_req(
        \request[3][0] ) );
  dccl_50 dccl_e ( .packet_addr_y_i({\packet_addr[1][3] , \packet_addr[1][2] , 
        \packet_addr[1][1] , \packet_addr[1][0] }), .packet_addr_x_i({
        \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] , 
        \packet_addr[1][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[1]), 
        .west_req(\request[2][1] ), .local_req(\request[3][1] ) );
  dccl_49 dccl_w ( .packet_addr_y_i({\packet_addr[2][3] , \packet_addr[2][2] , 
        \packet_addr[2][1] , \packet_addr[2][0] }), .packet_addr_x_i({
        \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] , 
        \packet_addr[2][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[2]), 
        .east_req(\request[1][1] ), .local_req(\request[3][2] ) );
  dccl_48 dccl_l ( .packet_addr_y_i({\packet_addr[3][3] , \packet_addr[3][2] , 
        \packet_addr[3][1] , \packet_addr[3][0] }), .packet_addr_x_i({
        \packet_addr[3][7] , \packet_addr[3][6] , \packet_addr[3][5] , 
        \packet_addr[3][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[3]), 
        .east_req(\request[1][2] ), .south_req(\request[0][0] ), .west_req(
        \request[2][2] ) );
endmodule


module mux3_1_19 ( data0, data1, data2, select0, select1, select2, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  output [15:0] data_o;
  input select0, select1, select2;
  wire   n1, n2, n6, n7, n8;

  AO222X1 U4 ( .IN1(data1[9]), .IN2(n8), .IN3(data0[9]), .IN4(n7), .IN5(
        data2[9]), .IN6(n6), .Q(data_o[9]) );
  AO222X1 U5 ( .IN1(data1[8]), .IN2(n8), .IN3(data0[8]), .IN4(n7), .IN5(
        data2[8]), .IN6(n6), .Q(data_o[8]) );
  AO222X1 U6 ( .IN1(data1[7]), .IN2(n8), .IN3(data0[7]), .IN4(n7), .IN5(
        data2[7]), .IN6(n6), .Q(data_o[7]) );
  AO222X1 U7 ( .IN1(data1[6]), .IN2(n8), .IN3(data0[6]), .IN4(n7), .IN5(
        data2[6]), .IN6(n6), .Q(data_o[6]) );
  AO222X1 U8 ( .IN1(data1[5]), .IN2(n8), .IN3(data0[5]), .IN4(n7), .IN5(
        data2[5]), .IN6(n6), .Q(data_o[5]) );
  AO222X1 U9 ( .IN1(data1[4]), .IN2(n8), .IN3(data0[4]), .IN4(n7), .IN5(
        data2[4]), .IN6(n6), .Q(data_o[4]) );
  AO222X1 U10 ( .IN1(data1[3]), .IN2(n8), .IN3(data0[3]), .IN4(n7), .IN5(
        data2[3]), .IN6(n6), .Q(data_o[3]) );
  AO222X1 U11 ( .IN1(data1[2]), .IN2(n8), .IN3(data0[2]), .IN4(n7), .IN5(
        data2[2]), .IN6(n6), .Q(data_o[2]) );
  AO222X1 U12 ( .IN1(data1[1]), .IN2(n8), .IN3(data0[1]), .IN4(n7), .IN5(
        data2[1]), .IN6(n6), .Q(data_o[1]) );
  AO222X1 U13 ( .IN1(data1[15]), .IN2(n8), .IN3(data0[15]), .IN4(n7), .IN5(
        data2[15]), .IN6(n6), .Q(data_o[15]) );
  AO222X1 U14 ( .IN1(data1[14]), .IN2(n8), .IN3(data0[14]), .IN4(n7), .IN5(
        data2[14]), .IN6(n6), .Q(data_o[14]) );
  AO222X1 U15 ( .IN1(data1[13]), .IN2(n8), .IN3(data0[13]), .IN4(n7), .IN5(
        data2[13]), .IN6(n6), .Q(data_o[13]) );
  AO222X1 U16 ( .IN1(data1[12]), .IN2(n8), .IN3(data0[12]), .IN4(n7), .IN5(
        data2[12]), .IN6(n6), .Q(data_o[12]) );
  AO222X1 U17 ( .IN1(data1[11]), .IN2(n8), .IN3(data0[11]), .IN4(n7), .IN5(
        data2[11]), .IN6(n6), .Q(data_o[11]) );
  AO222X1 U18 ( .IN1(data1[10]), .IN2(n8), .IN3(data0[10]), .IN4(n7), .IN5(
        data2[10]), .IN6(n6), .Q(data_o[10]) );
  AO222X1 U19 ( .IN1(data1[0]), .IN2(n8), .IN3(data0[0]), .IN4(n7), .IN5(
        data2[0]), .IN6(n6), .Q(data_o[0]) );
  INVX0 U2 ( .INP(select0), .ZN(n2) );
  INVX0 U3 ( .INP(select1), .ZN(n1) );
  AND3X1 U20 ( .IN1(n2), .IN2(n1), .IN3(select2), .Q(n6) );
  NOR3X0 U21 ( .IN1(select1), .IN2(select2), .IN3(n2), .QN(n7) );
  NOR3X0 U22 ( .IN1(select0), .IN2(select2), .IN3(n1), .QN(n8) );
endmodule


module mux3_1_18 ( data0, data1, data2, select0, select1, select2, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  output [15:0] data_o;
  input select0, select1, select2;
  wire   n1, n2, n6, n7, n8;

  AO222X1 U4 ( .IN1(data1[9]), .IN2(n8), .IN3(data0[9]), .IN4(n7), .IN5(
        data2[9]), .IN6(n6), .Q(data_o[9]) );
  AO222X1 U5 ( .IN1(data1[8]), .IN2(n8), .IN3(data0[8]), .IN4(n7), .IN5(
        data2[8]), .IN6(n6), .Q(data_o[8]) );
  AO222X1 U6 ( .IN1(data1[7]), .IN2(n8), .IN3(data0[7]), .IN4(n7), .IN5(
        data2[7]), .IN6(n6), .Q(data_o[7]) );
  AO222X1 U7 ( .IN1(data1[6]), .IN2(n8), .IN3(data0[6]), .IN4(n7), .IN5(
        data2[6]), .IN6(n6), .Q(data_o[6]) );
  AO222X1 U8 ( .IN1(data1[5]), .IN2(n8), .IN3(data0[5]), .IN4(n7), .IN5(
        data2[5]), .IN6(n6), .Q(data_o[5]) );
  AO222X1 U9 ( .IN1(data1[4]), .IN2(n8), .IN3(data0[4]), .IN4(n7), .IN5(
        data2[4]), .IN6(n6), .Q(data_o[4]) );
  AO222X1 U10 ( .IN1(data1[3]), .IN2(n8), .IN3(data0[3]), .IN4(n7), .IN5(
        data2[3]), .IN6(n6), .Q(data_o[3]) );
  AO222X1 U11 ( .IN1(data1[2]), .IN2(n8), .IN3(data0[2]), .IN4(n7), .IN5(
        data2[2]), .IN6(n6), .Q(data_o[2]) );
  AO222X1 U12 ( .IN1(data1[1]), .IN2(n8), .IN3(data0[1]), .IN4(n7), .IN5(
        data2[1]), .IN6(n6), .Q(data_o[1]) );
  AO222X1 U13 ( .IN1(data1[15]), .IN2(n8), .IN3(data0[15]), .IN4(n7), .IN5(
        data2[15]), .IN6(n6), .Q(data_o[15]) );
  AO222X1 U14 ( .IN1(data1[14]), .IN2(n8), .IN3(data0[14]), .IN4(n7), .IN5(
        data2[14]), .IN6(n6), .Q(data_o[14]) );
  AO222X1 U15 ( .IN1(data1[13]), .IN2(n8), .IN3(data0[13]), .IN4(n7), .IN5(
        data2[13]), .IN6(n6), .Q(data_o[13]) );
  AO222X1 U16 ( .IN1(data1[12]), .IN2(n8), .IN3(data0[12]), .IN4(n7), .IN5(
        data2[12]), .IN6(n6), .Q(data_o[12]) );
  AO222X1 U17 ( .IN1(data1[11]), .IN2(n8), .IN3(data0[11]), .IN4(n7), .IN5(
        data2[11]), .IN6(n6), .Q(data_o[11]) );
  AO222X1 U18 ( .IN1(data1[10]), .IN2(n8), .IN3(data0[10]), .IN4(n7), .IN5(
        data2[10]), .IN6(n6), .Q(data_o[10]) );
  AO222X1 U19 ( .IN1(data1[0]), .IN2(n8), .IN3(data0[0]), .IN4(n7), .IN5(
        data2[0]), .IN6(n6), .Q(data_o[0]) );
  INVX0 U2 ( .INP(select0), .ZN(n2) );
  INVX0 U3 ( .INP(select1), .ZN(n1) );
  AND3X1 U20 ( .IN1(n2), .IN2(n1), .IN3(select2), .Q(n6) );
  NOR3X0 U21 ( .IN1(select1), .IN2(select2), .IN3(n2), .QN(n7) );
  NOR3X0 U22 ( .IN1(select0), .IN2(select2), .IN3(n1), .QN(n8) );
endmodule


module mux3_1_17 ( data0, data1, data2, select0, select1, select2, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  output [15:0] data_o;
  input select0, select1, select2;
  wire   n1, n2, n6, n7, n8;

  AO222X1 U4 ( .IN1(data1[9]), .IN2(n8), .IN3(data0[9]), .IN4(n7), .IN5(
        data2[9]), .IN6(n6), .Q(data_o[9]) );
  AO222X1 U5 ( .IN1(data1[8]), .IN2(n8), .IN3(data0[8]), .IN4(n7), .IN5(
        data2[8]), .IN6(n6), .Q(data_o[8]) );
  AO222X1 U6 ( .IN1(data1[7]), .IN2(n8), .IN3(data0[7]), .IN4(n7), .IN5(
        data2[7]), .IN6(n6), .Q(data_o[7]) );
  AO222X1 U7 ( .IN1(data1[6]), .IN2(n8), .IN3(data0[6]), .IN4(n7), .IN5(
        data2[6]), .IN6(n6), .Q(data_o[6]) );
  AO222X1 U8 ( .IN1(data1[5]), .IN2(n8), .IN3(data0[5]), .IN4(n7), .IN5(
        data2[5]), .IN6(n6), .Q(data_o[5]) );
  AO222X1 U9 ( .IN1(data1[4]), .IN2(n8), .IN3(data0[4]), .IN4(n7), .IN5(
        data2[4]), .IN6(n6), .Q(data_o[4]) );
  AO222X1 U10 ( .IN1(data1[3]), .IN2(n8), .IN3(data0[3]), .IN4(n7), .IN5(
        data2[3]), .IN6(n6), .Q(data_o[3]) );
  AO222X1 U11 ( .IN1(data1[2]), .IN2(n8), .IN3(data0[2]), .IN4(n7), .IN5(
        data2[2]), .IN6(n6), .Q(data_o[2]) );
  AO222X1 U12 ( .IN1(data1[1]), .IN2(n8), .IN3(data0[1]), .IN4(n7), .IN5(
        data2[1]), .IN6(n6), .Q(data_o[1]) );
  AO222X1 U13 ( .IN1(data1[15]), .IN2(n8), .IN3(data0[15]), .IN4(n7), .IN5(
        data2[15]), .IN6(n6), .Q(data_o[15]) );
  AO222X1 U14 ( .IN1(data1[14]), .IN2(n8), .IN3(data0[14]), .IN4(n7), .IN5(
        data2[14]), .IN6(n6), .Q(data_o[14]) );
  AO222X1 U15 ( .IN1(data1[13]), .IN2(n8), .IN3(data0[13]), .IN4(n7), .IN5(
        data2[13]), .IN6(n6), .Q(data_o[13]) );
  AO222X1 U16 ( .IN1(data1[12]), .IN2(n8), .IN3(data0[12]), .IN4(n7), .IN5(
        data2[12]), .IN6(n6), .Q(data_o[12]) );
  AO222X1 U17 ( .IN1(data1[11]), .IN2(n8), .IN3(data0[11]), .IN4(n7), .IN5(
        data2[11]), .IN6(n6), .Q(data_o[11]) );
  AO222X1 U18 ( .IN1(data1[10]), .IN2(n8), .IN3(data0[10]), .IN4(n7), .IN5(
        data2[10]), .IN6(n6), .Q(data_o[10]) );
  AO222X1 U19 ( .IN1(data1[0]), .IN2(n8), .IN3(data0[0]), .IN4(n7), .IN5(
        data2[0]), .IN6(n6), .Q(data_o[0]) );
  INVX0 U2 ( .INP(select0), .ZN(n2) );
  INVX0 U3 ( .INP(select1), .ZN(n1) );
  AND3X1 U20 ( .IN1(n2), .IN2(n1), .IN3(select2), .Q(n6) );
  NOR3X0 U21 ( .IN1(select1), .IN2(select2), .IN3(n2), .QN(n7) );
  NOR3X0 U22 ( .IN1(select0), .IN2(select2), .IN3(n1), .QN(n8) );
endmodule



    module node4_NODE_X1_NODE_Y0I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__I_node_2_node_interface__ ( 
        \clk.clk , \reset.reset , \local_node.clk , 
        \local_node.buffer_full_in , \local_node.buffer_full_out , 
        \local_node.receiving_data , \local_node.sending_data , 
        \local_node.data_in , \local_node.data_out , \node_0.clk , 
        \node_0.buffer_full_in , \node_0.buffer_full_out , 
        \node_0.receiving_data , \node_0.sending_data , \node_0.data_in , 
        \node_0.data_out , \node_1.clk , \node_1.buffer_full_in , 
        \node_1.buffer_full_out , \node_1.receiving_data , 
        \node_1.sending_data , \node_1.data_in , \node_1.data_out , 
        \node_2.clk , \node_2.buffer_full_in , \node_2.buffer_full_out , 
        \node_2.receiving_data , \node_2.sending_data , \node_2.data_in , 
        \node_2.data_out  );
  input [15:0] \local_node.data_in ;
  output [15:0] \local_node.data_out ;
  input [15:0] \node_0.data_in ;
  output [15:0] \node_0.data_out ;
  input [15:0] \node_1.data_in ;
  output [15:0] \node_1.data_out ;
  input [15:0] \node_2.data_in ;
  output [15:0] \node_2.data_out ;
  input \clk.clk , \reset.reset , \local_node.buffer_full_in ,
         \local_node.receiving_data , \node_0.buffer_full_in ,
         \node_0.receiving_data , \node_1.buffer_full_in ,
         \node_1.receiving_data , \node_2.buffer_full_in ,
         \node_2.receiving_data ;
  output \local_node.buffer_full_out , \local_node.sending_data ,
         \node_0.buffer_full_out , \node_0.sending_data ,
         \node_1.buffer_full_out , \node_1.sending_data ,
         \node_2.buffer_full_out , \node_2.sending_data ;
  inout \local_node.clk ,  \node_0.clk ,  \node_1.clk ,  \node_2.clk ;
  wire   \buffer_out[3][15] , \buffer_out[3][14] , \buffer_out[3][13] ,
         \buffer_out[3][12] , \buffer_out[3][11] , \buffer_out[3][10] ,
         \buffer_out[3][9] , \buffer_out[3][8] , \buffer_out[3][7] ,
         \buffer_out[3][6] , \buffer_out[3][5] , \buffer_out[3][4] ,
         \buffer_out[3][3] , \buffer_out[3][2] , \buffer_out[3][1] ,
         \buffer_out[3][0] , \buffer_out[2][15] , \buffer_out[2][14] ,
         \buffer_out[2][13] , \buffer_out[2][12] , \buffer_out[2][11] ,
         \buffer_out[2][10] , \buffer_out[2][9] , \buffer_out[2][8] ,
         \buffer_out[2][7] , \buffer_out[2][6] , \buffer_out[2][5] ,
         \buffer_out[2][4] , \buffer_out[2][3] , \buffer_out[2][2] ,
         \buffer_out[2][1] , \buffer_out[2][0] , \buffer_out[1][15] ,
         \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] ,
         \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] ,
         \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] ,
         \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] ,
         \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] ,
         \buffer_out[0][15] , \buffer_out[0][14] , \buffer_out[0][13] ,
         \buffer_out[0][12] , \buffer_out[0][11] , \buffer_out[0][10] ,
         \buffer_out[0][9] , \buffer_out[0][8] , \buffer_out[0][7] ,
         \buffer_out[0][6] , \buffer_out[0][5] , \buffer_out[0][4] ,
         \buffer_out[0][3] , \buffer_out[0][2] , \buffer_out[0][1] ,
         \buffer_out[0][0] , \next_buffer_out[3][15] ,
         \next_buffer_out[3][14] , \next_buffer_out[3][13] ,
         \next_buffer_out[3][12] , \next_buffer_out[3][11] ,
         \next_buffer_out[3][10] , \next_buffer_out[3][9] ,
         \next_buffer_out[3][8] , \next_buffer_out[3][7] ,
         \next_buffer_out[3][6] , \next_buffer_out[3][5] ,
         \next_buffer_out[3][4] , \next_buffer_out[3][3] ,
         \next_buffer_out[3][2] , \next_buffer_out[3][1] ,
         \next_buffer_out[3][0] , \next_buffer_out[2][15] ,
         \next_buffer_out[2][14] , \next_buffer_out[2][13] ,
         \next_buffer_out[2][12] , \next_buffer_out[2][11] ,
         \next_buffer_out[2][10] , \next_buffer_out[2][9] ,
         \next_buffer_out[2][8] , \next_buffer_out[2][7] ,
         \next_buffer_out[2][6] , \next_buffer_out[2][5] ,
         \next_buffer_out[2][4] , \next_buffer_out[2][3] ,
         \next_buffer_out[2][2] , \next_buffer_out[2][1] ,
         \next_buffer_out[2][0] , \next_buffer_out[1][15] ,
         \next_buffer_out[1][14] , \next_buffer_out[1][13] ,
         \next_buffer_out[1][12] , \next_buffer_out[1][11] ,
         \next_buffer_out[1][10] , \next_buffer_out[1][9] ,
         \next_buffer_out[1][8] , \next_buffer_out[1][7] ,
         \next_buffer_out[1][6] , \next_buffer_out[1][5] ,
         \next_buffer_out[1][4] , \next_buffer_out[1][3] ,
         \next_buffer_out[1][2] , \next_buffer_out[1][1] ,
         \next_buffer_out[1][0] , \next_buffer_out[0][15] ,
         \next_buffer_out[0][14] , \next_buffer_out[0][13] ,
         \next_buffer_out[0][12] , \next_buffer_out[0][11] ,
         \next_buffer_out[0][10] , \next_buffer_out[0][9] ,
         \next_buffer_out[0][8] , \next_buffer_out[0][7] ,
         \next_buffer_out[0][6] , \next_buffer_out[0][5] ,
         \next_buffer_out[0][4] , \next_buffer_out[0][3] ,
         \next_buffer_out[0][2] , \next_buffer_out[0][1] ,
         \next_buffer_out[0][0] ;
  wire   [3:0] buffer_full_in;
  wire   [3:0] receiving_data;
  wire   [3:0] pop_v;
  wire   [3:0] data_valid;
  wire   [3:0] next_data_valid;
  wire   [2:0] grant_1;
  wire   [2:0] grant_2;
  wire   [2:0] grant_3;
  tri   \local_node.buffer_full_in ;
  tri   \local_node.buffer_full_out ;
  tri   \local_node.receiving_data ;
  tri   \local_node.sending_data ;
  tri   [15:0] \local_node.data_in ;
  tri   [15:0] \local_node.data_out ;

  converter_out_I_n_node_interface_dut_ c3 ( .\n.buffer_full_in (
        \local_node.buffer_full_in ), .\n.receiving_data (
        \local_node.receiving_data ), .\n.data_in (\local_node.data_in ), 
        .\n.buffer_full_out (\local_node.buffer_full_out ), .\n.sending_data (
        \local_node.sending_data ), .\n.data_out (\local_node.data_out ), 
        .buffer_full_in(1'b0), .receiving_data(1'b0), .data_in({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  fifo_kev_51 \genblk1[0].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[0]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[0]), .data_out({\buffer_out[0][15] , 
        \buffer_out[0][14] , \buffer_out[0][13] , \buffer_out[0][12] , 
        \buffer_out[0][11] , \buffer_out[0][10] , \buffer_out[0][9] , 
        \buffer_out[0][8] , \buffer_out[0][7] , \buffer_out[0][6] , 
        \buffer_out[0][5] , \buffer_out[0][4] , \buffer_out[0][3] , 
        \buffer_out[0][2] , \buffer_out[0][1] , \buffer_out[0][0] }), 
        .next_data_out({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] , 
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .next_data_valid(
        next_data_valid[0]) );
  address_counter_51 \genblk1[0].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] }), 
        .buffer_data_valid(next_data_valid[0]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .buffer_pop(
        pop_v[0]), .receiving_data(1'b0) );
  fifo_kev_50 \genblk1[1].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[1]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[1]), .data_out({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), 
        .next_data_out({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] , 
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .next_data_valid(
        next_data_valid[1]) );
  address_counter_50 \genblk1[1].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] }), 
        .buffer_data_valid(next_data_valid[1]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .buffer_pop(
        pop_v[1]), .receiving_data(1'b0) );
  fifo_kev_49 \genblk1[2].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[2]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[2]), .data_out({\buffer_out[2][15] , 
        \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] , 
        \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] , 
        \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] , 
        \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] , 
        \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] }), 
        .next_data_out({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] , 
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .next_data_valid(
        next_data_valid[2]) );
  address_counter_49 \genblk1[2].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] }), 
        .buffer_data_valid(next_data_valid[2]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .buffer_pop(
        pop_v[2]), .receiving_data(1'b0) );
  fifo_kev_48 \genblk1[3].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[3]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[3]), .data_out({\buffer_out[3][15] , 
        \buffer_out[3][14] , \buffer_out[3][13] , \buffer_out[3][12] , 
        \buffer_out[3][11] , \buffer_out[3][10] , \buffer_out[3][9] , 
        \buffer_out[3][8] , \buffer_out[3][7] , \buffer_out[3][6] , 
        \buffer_out[3][5] , \buffer_out[3][4] , \buffer_out[3][3] , 
        \buffer_out[3][2] , \buffer_out[3][1] , \buffer_out[3][0] }), 
        .next_data_out({\next_buffer_out[3][15] , \next_buffer_out[3][14] , 
        \next_buffer_out[3][13] , \next_buffer_out[3][12] , 
        \next_buffer_out[3][11] , \next_buffer_out[3][10] , 
        \next_buffer_out[3][9] , \next_buffer_out[3][8] , 
        \next_buffer_out[3][7] , \next_buffer_out[3][6] , 
        \next_buffer_out[3][5] , \next_buffer_out[3][4] , 
        \next_buffer_out[3][3] , \next_buffer_out[3][2] , 
        \next_buffer_out[3][1] , \next_buffer_out[3][0] }), .next_data_valid(
        next_data_valid[3]) );
  address_counter_48 \genblk1[3].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[3][15] , \next_buffer_out[3][14] , 
        \next_buffer_out[3][13] , \next_buffer_out[3][12] , 
        \next_buffer_out[3][11] , \next_buffer_out[3][10] , 
        \next_buffer_out[3][9] , \next_buffer_out[3][8] }), 
        .buffer_data_valid(next_data_valid[3]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[3][7] , \next_buffer_out[3][6] , 
        \next_buffer_out[3][5] , \next_buffer_out[3][4] , 
        \next_buffer_out[3][3] , \next_buffer_out[3][2] , 
        \next_buffer_out[3][1] , \next_buffer_out[3][0] }), .buffer_pop(
        pop_v[3]), .receiving_data(1'b0) );
  converter_out_I_n_node_interface_dut_ \genblk2.c0  ( .\n.buffer_full_in (
        \node_0.buffer_full_in ), .\n.receiving_data (\node_0.receiving_data ), 
        .\n.data_in (\node_0.data_in ), .\n.buffer_full_out (
        \node_0.buffer_full_out ), .\n.sending_data (\node_0.sending_data ), 
        .\n.data_out (\node_0.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_in_I_n_node_interface_dut__19 \genblk2.c1  ( .\n.buffer_full_in (
        \node_1.buffer_full_in ), .\n.receiving_data (\node_1.receiving_data ), 
        .\n.data_in (\node_1.data_in ), .\n.buffer_full_out (
        \node_1.buffer_full_out ), .\n.sending_data (\node_1.sending_data ), 
        .\n.data_out (\node_1.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_out_I_n_node_interface_dut_ \genblk2.c2  ( .\n.buffer_full_in (
        \node_2.buffer_full_in ), .\n.receiving_data (\node_2.receiving_data ), 
        .\n.data_in (\node_2.data_in ), .\n.buffer_full_out (
        \node_2.buffer_full_out ), .\n.sending_data (\node_2.sending_data ), 
        .\n.data_out (\node_2.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  controller4_edge_n_1 \genblk2.n  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .packet_addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .local_addr({1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .packet_valid(data_valid), .buffer_full_in({1'b0, 1'b0, 1'b0, 1'b0}), 
        .grant_1(grant_1), .grant_2(grant_2), .grant_3(grant_3), .pop_v(pop_v)
         );
  mux3_1_19 \genblk2.mux_e  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[2][15] , 
        \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] , 
        \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] , 
        \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] , 
        \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] , 
        \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] }), .data2({
        \buffer_out[3][15] , \buffer_out[3][14] , \buffer_out[3][13] , 
        \buffer_out[3][12] , \buffer_out[3][11] , \buffer_out[3][10] , 
        \buffer_out[3][9] , \buffer_out[3][8] , \buffer_out[3][7] , 
        \buffer_out[3][6] , \buffer_out[3][5] , \buffer_out[3][4] , 
        \buffer_out[3][3] , \buffer_out[3][2] , \buffer_out[3][1] , 
        \buffer_out[3][0] }), .select0(grant_1[0]), .select1(grant_1[1]), 
        .select2(grant_1[2]) );
  mux3_1_18 \genblk2.mux_w  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[3][15] , \buffer_out[3][14] , \buffer_out[3][13] , 
        \buffer_out[3][12] , \buffer_out[3][11] , \buffer_out[3][10] , 
        \buffer_out[3][9] , \buffer_out[3][8] , \buffer_out[3][7] , 
        \buffer_out[3][6] , \buffer_out[3][5] , \buffer_out[3][4] , 
        \buffer_out[3][3] , \buffer_out[3][2] , \buffer_out[3][1] , 
        \buffer_out[3][0] }), .select0(grant_2[0]), .select1(grant_2[1]), 
        .select2(grant_2[2]) );
  mux3_1_17 \genblk2.mux_l  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[2][15] , \buffer_out[2][14] , \buffer_out[2][13] , 
        \buffer_out[2][12] , \buffer_out[2][11] , \buffer_out[2][10] , 
        \buffer_out[2][9] , \buffer_out[2][8] , \buffer_out[2][7] , 
        \buffer_out[2][6] , \buffer_out[2][5] , \buffer_out[2][4] , 
        \buffer_out[2][3] , \buffer_out[2][2] , \buffer_out[2][1] , 
        \buffer_out[2][0] }), .select0(grant_3[0]), .select1(grant_3[1]), 
        .select2(grant_3[2]) );
endmodule


module fifo_kev_47 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_95 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_47 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_95 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_94 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_47 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_94 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_47_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_47 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_47 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_47 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_47_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_46 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_93 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_46 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_93 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_92 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_46 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_92 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_46_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_46 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_46 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_46 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_46_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_45 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_91 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_45 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_91 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_90 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_45 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_90 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_45_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_45 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_45 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_45 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_45_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_44 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_89 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_44 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_89 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_88 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_44 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_88 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_44_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_44 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_44 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_44 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_44_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module converter_in_I_n_node_interface_dut__18 ( \n.buffer_full_in , 
        \n.receiving_data , \n.data_in , \n.buffer_full_out , \n.sending_data , 
        \n.data_out , buffer_full_out, sending_data, data_out, buffer_full_in, 
        receiving_data, data_in );
  input [15:0] \n.data_in ;
  output [15:0] \n.data_out ;
  output [15:0] data_out;
  input [15:0] data_in;
  input \n.buffer_full_in , \n.receiving_data , buffer_full_in, receiving_data;
  output \n.buffer_full_out , \n.sending_data , buffer_full_out, sending_data;
  wire   \n.buffer_full_in , \n.receiving_data , buffer_full_in,
         receiving_data;
  assign buffer_full_out = \n.buffer_full_in ;
  assign sending_data = \n.receiving_data ;
  assign data_out[15] = \n.data_in  [15];
  assign data_out[14] = \n.data_in  [14];
  assign data_out[13] = \n.data_in  [13];
  assign data_out[12] = \n.data_in  [12];
  assign data_out[11] = \n.data_in  [11];
  assign data_out[10] = \n.data_in  [10];
  assign data_out[9] = \n.data_in  [9];
  assign data_out[8] = \n.data_in  [8];
  assign data_out[7] = \n.data_in  [7];
  assign data_out[6] = \n.data_in  [6];
  assign data_out[5] = \n.data_in  [5];
  assign data_out[4] = \n.data_in  [4];
  assign data_out[3] = \n.data_in  [3];
  assign data_out[2] = \n.data_in  [2];
  assign data_out[1] = \n.data_in  [1];
  assign data_out[0] = \n.data_in  [0];
  assign \n.buffer_full_out  = buffer_full_in;
  assign \n.sending_data  = receiving_data;
  assign \n.data_out  [15] = data_in[15];
  assign \n.data_out  [14] = data_in[14];
  assign \n.data_out  [13] = data_in[13];
  assign \n.data_out  [12] = data_in[12];
  assign \n.data_out  [11] = data_in[11];
  assign \n.data_out  [10] = data_in[10];
  assign \n.data_out  [9] = data_in[9];
  assign \n.data_out  [8] = data_in[8];
  assign \n.data_out  [7] = data_in[7];
  assign \n.data_out  [6] = data_in[6];
  assign \n.data_out  [5] = data_in[5];
  assign \n.data_out  [4] = data_in[4];
  assign \n.data_out  [3] = data_in[3];
  assign \n.data_out  [2] = data_in[2];
  assign \n.data_out  [1] = data_in[1];
  assign \n.data_out  [0] = data_in[0];

endmodule


module flipflop_BITS3_33 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_33 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_33 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS3_32 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_32 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_32 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS1_73 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_73 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_73 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_72 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_72 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_72 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter3_16 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [2:0] request;
  output [2:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[1][2] , \req_i[1][1] , \req_i[1][0] , \req_i[0][2] ,
         \req_i[0][1] , tail_en, N99, N100, N101, N110, N111, N118, N119, N120,
         N121, n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [1:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N99 = request[0];
  assign N100 = request[1];
  assign N101 = request[2];

  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(N111), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(N110), .Q(\req_i[0][1] ) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N121), .D(tail_en), .Q(req_en[0]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N120), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N119), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N118), .Q(grant[0]) );
  AND2X1 U20 ( .IN1(n8), .IN2(N101), .Q(n7) );
  OR3X1 U21 ( .IN1(n3), .IN2(N111), .IN3(n6), .Q(N121) );
  NOR3X0 U22 ( .IN1(N99), .IN2(N100), .IN3(n6), .QN(N120) );
  NOR3X0 U23 ( .IN1(n2), .IN2(N99), .IN3(n6), .QN(N119) );
  NAND3X0 U24 ( .IN1(n2), .IN2(n3), .IN3(n1), .QN(n5) );
  AO22X1 U25 ( .IN1(N100), .IN2(N101), .IN3(N99), .IN4(N101), .Q(N111) );
  INVX0 U10 ( .INP(N101), .ZN(n3) );
  NAND2X1 U11 ( .IN1(n5), .IN2(n4), .QN(n6) );
  INVX0 U12 ( .INP(N99), .ZN(n1) );
  INVX0 U13 ( .INP(N100), .ZN(n2) );
  INVX0 U14 ( .INP(buffer_full_i), .ZN(n4) );
  NAND2X1 U15 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NOR2X0 U16 ( .IN1(n1), .IN2(n6), .QN(N118) );
  NOR2X0 U17 ( .IN1(n1), .IN2(n2), .QN(N110) );
  OA21X1 U18 ( .IN1(N110), .IN2(n7), .IN3(n4), .Q(tail_en) );
  OA21X1 U19 ( .IN1(N101), .IN2(n8), .IN3(n4), .Q(grant_v_o) );
  register_BITS3_33 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][2] , \req_i[0][1] , 1'b0}), .data_o({
        1'b0, 1'b0, 1'b0}) );
  register_BITS3_32 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][2] , \req_i[1][1] , \req_i[1][0] }), 
        .data_o({1'b0, 1'b0, 1'b0}) );
  register_BITS1_73 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b1), .data_o(1'b0) );
  register_BITS1_72 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module flipflop_BITS3_31 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_31 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_31 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS3_30 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_30 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_30 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS1_71 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_71 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_71 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_70 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_70 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_70 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter3_15 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [2:0] request;
  output [2:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[1][2] , \req_i[1][1] , \req_i[1][0] , \req_i[0][2] ,
         \req_i[0][1] , tail_en, N99, N100, N101, N110, N111, N118, N119, N120,
         N121, n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [1:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N99 = request[0];
  assign N100 = request[1];
  assign N101 = request[2];

  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(N111), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(N110), .Q(\req_i[0][1] ) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N121), .D(tail_en), .Q(req_en[0]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N120), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N119), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N118), .Q(grant[0]) );
  AND2X1 U20 ( .IN1(n8), .IN2(N101), .Q(n7) );
  OR3X1 U21 ( .IN1(n3), .IN2(N111), .IN3(n6), .Q(N121) );
  NOR3X0 U22 ( .IN1(N99), .IN2(N100), .IN3(n6), .QN(N120) );
  NOR3X0 U23 ( .IN1(n2), .IN2(N99), .IN3(n6), .QN(N119) );
  NAND3X0 U24 ( .IN1(n2), .IN2(n3), .IN3(n1), .QN(n5) );
  AO22X1 U25 ( .IN1(N100), .IN2(N101), .IN3(N99), .IN4(N101), .Q(N111) );
  INVX0 U10 ( .INP(N101), .ZN(n3) );
  NAND2X1 U11 ( .IN1(n5), .IN2(n4), .QN(n6) );
  INVX0 U12 ( .INP(N99), .ZN(n1) );
  INVX0 U13 ( .INP(N100), .ZN(n2) );
  INVX0 U14 ( .INP(buffer_full_i), .ZN(n4) );
  NAND2X1 U15 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NOR2X0 U16 ( .IN1(n1), .IN2(n6), .QN(N118) );
  NOR2X0 U17 ( .IN1(n1), .IN2(n2), .QN(N110) );
  OA21X1 U18 ( .IN1(N110), .IN2(n7), .IN3(n4), .Q(tail_en) );
  OA21X1 U19 ( .IN1(N101), .IN2(n8), .IN3(n4), .Q(grant_v_o) );
  register_BITS3_31 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][2] , \req_i[0][1] , 1'b0}), .data_o({
        1'b0, 1'b0, 1'b0}) );
  register_BITS3_30 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][2] , \req_i[1][1] , \req_i[1][0] }), 
        .data_o({1'b0, 1'b0, 1'b0}) );
  register_BITS1_71 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b1), .data_o(1'b0) );
  register_BITS1_70 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module flipflop_BITS3_29 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_29 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_29 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS3_28 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_28 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_28 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS1_69 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_69 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_69 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_68 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_68 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_68 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter3_14 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [2:0] request;
  output [2:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[1][2] , \req_i[1][1] , \req_i[1][0] , \req_i[0][2] ,
         \req_i[0][1] , tail_en, N99, N100, N101, N110, N111, N118, N119, N120,
         N121, n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [1:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N99 = request[0];
  assign N100 = request[1];
  assign N101 = request[2];

  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(N111), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(N110), .Q(\req_i[0][1] ) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N121), .D(tail_en), .Q(req_en[0]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N120), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N119), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N118), .Q(grant[0]) );
  AND2X1 U20 ( .IN1(n8), .IN2(N101), .Q(n7) );
  OR3X1 U21 ( .IN1(n3), .IN2(N111), .IN3(n6), .Q(N121) );
  NOR3X0 U22 ( .IN1(N99), .IN2(N100), .IN3(n6), .QN(N120) );
  NOR3X0 U23 ( .IN1(n2), .IN2(N99), .IN3(n6), .QN(N119) );
  NAND3X0 U24 ( .IN1(n2), .IN2(n3), .IN3(n1), .QN(n5) );
  AO22X1 U25 ( .IN1(N100), .IN2(N101), .IN3(N99), .IN4(N101), .Q(N111) );
  INVX0 U10 ( .INP(N101), .ZN(n3) );
  NAND2X1 U11 ( .IN1(n5), .IN2(n4), .QN(n6) );
  INVX0 U12 ( .INP(N99), .ZN(n1) );
  INVX0 U13 ( .INP(N100), .ZN(n2) );
  INVX0 U14 ( .INP(buffer_full_i), .ZN(n4) );
  NAND2X1 U15 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NOR2X0 U16 ( .IN1(n1), .IN2(n6), .QN(N118) );
  NOR2X0 U17 ( .IN1(n1), .IN2(n2), .QN(N110) );
  OA21X1 U18 ( .IN1(N110), .IN2(n7), .IN3(n4), .Q(tail_en) );
  OA21X1 U19 ( .IN1(N101), .IN2(n8), .IN3(n4), .Q(grant_v_o) );
  register_BITS3_29 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][2] , \req_i[0][1] , 1'b0}), .data_o({
        1'b0, 1'b0, 1'b0}) );
  register_BITS3_28 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][2] , \req_i[1][1] , \req_i[1][0] }), 
        .data_o({1'b0, 1'b0, 1'b0}) );
  register_BITS1_69 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b1), .data_o(1'b0) );
  register_BITS1_68 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module dccl_47 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_46 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_45 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_44 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module controller4_edge_n_0 ( clk, rst, .packet_addr({\packet_addr[3][7] , 
        \packet_addr[3][6] , \packet_addr[3][5] , \packet_addr[3][4] , 
        \packet_addr[3][3] , \packet_addr[3][2] , \packet_addr[3][1] , 
        \packet_addr[3][0] , \packet_addr[2][7] , \packet_addr[2][6] , 
        \packet_addr[2][5] , \packet_addr[2][4] , \packet_addr[2][3] , 
        \packet_addr[2][2] , \packet_addr[2][1] , \packet_addr[2][0] , 
        \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] , 
        \packet_addr[1][4] , \packet_addr[1][3] , \packet_addr[1][2] , 
        \packet_addr[1][1] , \packet_addr[1][0] , \packet_addr[0][7] , 
        \packet_addr[0][6] , \packet_addr[0][5] , \packet_addr[0][4] , 
        \packet_addr[0][3] , \packet_addr[0][2] , \packet_addr[0][1] , 
        \packet_addr[0][0] }), local_addr, packet_valid, buffer_full_in, 
        grant_1, grant_2, grant_3, grant_v, pop_v );
  input [7:0] local_addr;
  input [3:0] packet_valid;
  input [3:0] buffer_full_in;
  output [2:0] grant_1;
  output [2:0] grant_2;
  output [2:0] grant_3;
  output [3:0] grant_v;
  output [3:0] pop_v;
  input clk, rst, \packet_addr[3][7] , \packet_addr[3][6] ,
         \packet_addr[3][5] , \packet_addr[3][4] , \packet_addr[3][3] ,
         \packet_addr[3][2] , \packet_addr[3][1] , \packet_addr[3][0] ,
         \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] ,
         \packet_addr[2][4] , \packet_addr[2][3] , \packet_addr[2][2] ,
         \packet_addr[2][1] , \packet_addr[2][0] , \packet_addr[1][7] ,
         \packet_addr[1][6] , \packet_addr[1][5] , \packet_addr[1][4] ,
         \packet_addr[1][3] , \packet_addr[1][2] , \packet_addr[1][1] ,
         \packet_addr[1][0] , \packet_addr[0][7] , \packet_addr[0][6] ,
         \packet_addr[0][5] , \packet_addr[0][4] , \packet_addr[0][3] ,
         \packet_addr[0][2] , \packet_addr[0][1] , \packet_addr[0][0] ;
  wire   \request[3][2] , \request[3][1] , \request[3][0] , \request[2][2] ,
         \request[2][1] , \request[2][0] , \request[1][2] , \request[1][1] ,
         \request[1][0] , \request[0][0] , n1;

  OR3X1 U3 ( .IN1(grant_2[2]), .IN2(grant_1[2]), .IN3(grant_v[0]), .Q(pop_v[3]) );
  OR2X1 U4 ( .IN1(grant_1[1]), .IN2(grant_3[2]), .Q(pop_v[2]) );
  OR2X1 U5 ( .IN1(grant_2[1]), .IN2(grant_3[1]), .Q(pop_v[1]) );
  OR3X1 U6 ( .IN1(grant_3[0]), .IN2(grant_2[0]), .IN3(grant_1[0]), .Q(pop_v[0]) );
  NOR2X0 U1 ( .IN1(n1), .IN2(buffer_full_in[0]), .QN(grant_v[0]) );
  INVX0 U2 ( .INP(\request[0][0] ), .ZN(n1) );
  arbiter3_16 arbiter_e ( .clk(clk), .rst(rst), .request({\request[1][2] , 
        \request[1][1] , \request[1][0] }), .buffer_full_i(buffer_full_in[1]), 
        .grant(grant_1), .grant_v_o(grant_v[1]) );
  arbiter3_15 arbiter_w ( .clk(clk), .rst(rst), .request({\request[2][2] , 
        \request[2][1] , \request[2][0] }), .buffer_full_i(buffer_full_in[2]), 
        .grant(grant_2), .grant_v_o(grant_v[2]) );
  arbiter3_14 arbiter_l ( .clk(clk), .rst(rst), .request({\request[3][2] , 
        \request[3][1] , \request[3][0] }), .buffer_full_i(buffer_full_in[3]), 
        .grant(grant_3), .grant_v_o(grant_v[3]) );
  dccl_47 dccl_s ( .packet_addr_y_i({\packet_addr[0][3] , \packet_addr[0][2] , 
        \packet_addr[0][1] , \packet_addr[0][0] }), .packet_addr_x_i({
        \packet_addr[0][7] , \packet_addr[0][6] , \packet_addr[0][5] , 
        \packet_addr[0][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[0]), 
        .east_req(\request[1][0] ), .west_req(\request[2][0] ), .local_req(
        \request[3][0] ) );
  dccl_46 dccl_e ( .packet_addr_y_i({\packet_addr[1][3] , \packet_addr[1][2] , 
        \packet_addr[1][1] , \packet_addr[1][0] }), .packet_addr_x_i({
        \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] , 
        \packet_addr[1][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[1]), 
        .west_req(\request[2][1] ), .local_req(\request[3][1] ) );
  dccl_45 dccl_w ( .packet_addr_y_i({\packet_addr[2][3] , \packet_addr[2][2] , 
        \packet_addr[2][1] , \packet_addr[2][0] }), .packet_addr_x_i({
        \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] , 
        \packet_addr[2][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[2]), 
        .east_req(\request[1][1] ), .local_req(\request[3][2] ) );
  dccl_44 dccl_l ( .packet_addr_y_i({\packet_addr[3][3] , \packet_addr[3][2] , 
        \packet_addr[3][1] , \packet_addr[3][0] }), .packet_addr_x_i({
        \packet_addr[3][7] , \packet_addr[3][6] , \packet_addr[3][5] , 
        \packet_addr[3][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[3]), 
        .east_req(\request[1][2] ), .south_req(\request[0][0] ), .west_req(
        \request[2][2] ) );
endmodule


module mux3_1_16 ( data0, data1, data2, select0, select1, select2, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  output [15:0] data_o;
  input select0, select1, select2;
  wire   n1, n2, n6, n7, n8;

  AO222X1 U4 ( .IN1(data1[9]), .IN2(n8), .IN3(data0[9]), .IN4(n7), .IN5(
        data2[9]), .IN6(n6), .Q(data_o[9]) );
  AO222X1 U5 ( .IN1(data1[8]), .IN2(n8), .IN3(data0[8]), .IN4(n7), .IN5(
        data2[8]), .IN6(n6), .Q(data_o[8]) );
  AO222X1 U6 ( .IN1(data1[7]), .IN2(n8), .IN3(data0[7]), .IN4(n7), .IN5(
        data2[7]), .IN6(n6), .Q(data_o[7]) );
  AO222X1 U7 ( .IN1(data1[6]), .IN2(n8), .IN3(data0[6]), .IN4(n7), .IN5(
        data2[6]), .IN6(n6), .Q(data_o[6]) );
  AO222X1 U8 ( .IN1(data1[5]), .IN2(n8), .IN3(data0[5]), .IN4(n7), .IN5(
        data2[5]), .IN6(n6), .Q(data_o[5]) );
  AO222X1 U9 ( .IN1(data1[4]), .IN2(n8), .IN3(data0[4]), .IN4(n7), .IN5(
        data2[4]), .IN6(n6), .Q(data_o[4]) );
  AO222X1 U10 ( .IN1(data1[3]), .IN2(n8), .IN3(data0[3]), .IN4(n7), .IN5(
        data2[3]), .IN6(n6), .Q(data_o[3]) );
  AO222X1 U11 ( .IN1(data1[2]), .IN2(n8), .IN3(data0[2]), .IN4(n7), .IN5(
        data2[2]), .IN6(n6), .Q(data_o[2]) );
  AO222X1 U12 ( .IN1(data1[1]), .IN2(n8), .IN3(data0[1]), .IN4(n7), .IN5(
        data2[1]), .IN6(n6), .Q(data_o[1]) );
  AO222X1 U13 ( .IN1(data1[15]), .IN2(n8), .IN3(data0[15]), .IN4(n7), .IN5(
        data2[15]), .IN6(n6), .Q(data_o[15]) );
  AO222X1 U14 ( .IN1(data1[14]), .IN2(n8), .IN3(data0[14]), .IN4(n7), .IN5(
        data2[14]), .IN6(n6), .Q(data_o[14]) );
  AO222X1 U15 ( .IN1(data1[13]), .IN2(n8), .IN3(data0[13]), .IN4(n7), .IN5(
        data2[13]), .IN6(n6), .Q(data_o[13]) );
  AO222X1 U16 ( .IN1(data1[12]), .IN2(n8), .IN3(data0[12]), .IN4(n7), .IN5(
        data2[12]), .IN6(n6), .Q(data_o[12]) );
  AO222X1 U17 ( .IN1(data1[11]), .IN2(n8), .IN3(data0[11]), .IN4(n7), .IN5(
        data2[11]), .IN6(n6), .Q(data_o[11]) );
  AO222X1 U18 ( .IN1(data1[10]), .IN2(n8), .IN3(data0[10]), .IN4(n7), .IN5(
        data2[10]), .IN6(n6), .Q(data_o[10]) );
  AO222X1 U19 ( .IN1(data1[0]), .IN2(n8), .IN3(data0[0]), .IN4(n7), .IN5(
        data2[0]), .IN6(n6), .Q(data_o[0]) );
  INVX0 U2 ( .INP(select0), .ZN(n2) );
  INVX0 U3 ( .INP(select1), .ZN(n1) );
  AND3X1 U20 ( .IN1(n2), .IN2(n1), .IN3(select2), .Q(n6) );
  NOR3X0 U21 ( .IN1(select1), .IN2(select2), .IN3(n2), .QN(n7) );
  NOR3X0 U22 ( .IN1(select0), .IN2(select2), .IN3(n1), .QN(n8) );
endmodule


module mux3_1_15 ( data0, data1, data2, select0, select1, select2, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  output [15:0] data_o;
  input select0, select1, select2;
  wire   n1, n2, n6, n7, n8;

  AO222X1 U4 ( .IN1(data1[9]), .IN2(n8), .IN3(data0[9]), .IN4(n7), .IN5(
        data2[9]), .IN6(n6), .Q(data_o[9]) );
  AO222X1 U5 ( .IN1(data1[8]), .IN2(n8), .IN3(data0[8]), .IN4(n7), .IN5(
        data2[8]), .IN6(n6), .Q(data_o[8]) );
  AO222X1 U6 ( .IN1(data1[7]), .IN2(n8), .IN3(data0[7]), .IN4(n7), .IN5(
        data2[7]), .IN6(n6), .Q(data_o[7]) );
  AO222X1 U7 ( .IN1(data1[6]), .IN2(n8), .IN3(data0[6]), .IN4(n7), .IN5(
        data2[6]), .IN6(n6), .Q(data_o[6]) );
  AO222X1 U8 ( .IN1(data1[5]), .IN2(n8), .IN3(data0[5]), .IN4(n7), .IN5(
        data2[5]), .IN6(n6), .Q(data_o[5]) );
  AO222X1 U9 ( .IN1(data1[4]), .IN2(n8), .IN3(data0[4]), .IN4(n7), .IN5(
        data2[4]), .IN6(n6), .Q(data_o[4]) );
  AO222X1 U10 ( .IN1(data1[3]), .IN2(n8), .IN3(data0[3]), .IN4(n7), .IN5(
        data2[3]), .IN6(n6), .Q(data_o[3]) );
  AO222X1 U11 ( .IN1(data1[2]), .IN2(n8), .IN3(data0[2]), .IN4(n7), .IN5(
        data2[2]), .IN6(n6), .Q(data_o[2]) );
  AO222X1 U12 ( .IN1(data1[1]), .IN2(n8), .IN3(data0[1]), .IN4(n7), .IN5(
        data2[1]), .IN6(n6), .Q(data_o[1]) );
  AO222X1 U13 ( .IN1(data1[15]), .IN2(n8), .IN3(data0[15]), .IN4(n7), .IN5(
        data2[15]), .IN6(n6), .Q(data_o[15]) );
  AO222X1 U14 ( .IN1(data1[14]), .IN2(n8), .IN3(data0[14]), .IN4(n7), .IN5(
        data2[14]), .IN6(n6), .Q(data_o[14]) );
  AO222X1 U15 ( .IN1(data1[13]), .IN2(n8), .IN3(data0[13]), .IN4(n7), .IN5(
        data2[13]), .IN6(n6), .Q(data_o[13]) );
  AO222X1 U16 ( .IN1(data1[12]), .IN2(n8), .IN3(data0[12]), .IN4(n7), .IN5(
        data2[12]), .IN6(n6), .Q(data_o[12]) );
  AO222X1 U17 ( .IN1(data1[11]), .IN2(n8), .IN3(data0[11]), .IN4(n7), .IN5(
        data2[11]), .IN6(n6), .Q(data_o[11]) );
  AO222X1 U18 ( .IN1(data1[10]), .IN2(n8), .IN3(data0[10]), .IN4(n7), .IN5(
        data2[10]), .IN6(n6), .Q(data_o[10]) );
  AO222X1 U19 ( .IN1(data1[0]), .IN2(n8), .IN3(data0[0]), .IN4(n7), .IN5(
        data2[0]), .IN6(n6), .Q(data_o[0]) );
  INVX0 U2 ( .INP(select0), .ZN(n2) );
  INVX0 U3 ( .INP(select1), .ZN(n1) );
  AND3X1 U20 ( .IN1(n2), .IN2(n1), .IN3(select2), .Q(n6) );
  NOR3X0 U21 ( .IN1(select1), .IN2(select2), .IN3(n2), .QN(n7) );
  NOR3X0 U22 ( .IN1(select0), .IN2(select2), .IN3(n1), .QN(n8) );
endmodule


module mux3_1_14 ( data0, data1, data2, select0, select1, select2, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  output [15:0] data_o;
  input select0, select1, select2;
  wire   n1, n2, n6, n7, n8;

  AO222X1 U4 ( .IN1(data1[9]), .IN2(n8), .IN3(data0[9]), .IN4(n7), .IN5(
        data2[9]), .IN6(n6), .Q(data_o[9]) );
  AO222X1 U5 ( .IN1(data1[8]), .IN2(n8), .IN3(data0[8]), .IN4(n7), .IN5(
        data2[8]), .IN6(n6), .Q(data_o[8]) );
  AO222X1 U6 ( .IN1(data1[7]), .IN2(n8), .IN3(data0[7]), .IN4(n7), .IN5(
        data2[7]), .IN6(n6), .Q(data_o[7]) );
  AO222X1 U7 ( .IN1(data1[6]), .IN2(n8), .IN3(data0[6]), .IN4(n7), .IN5(
        data2[6]), .IN6(n6), .Q(data_o[6]) );
  AO222X1 U8 ( .IN1(data1[5]), .IN2(n8), .IN3(data0[5]), .IN4(n7), .IN5(
        data2[5]), .IN6(n6), .Q(data_o[5]) );
  AO222X1 U9 ( .IN1(data1[4]), .IN2(n8), .IN3(data0[4]), .IN4(n7), .IN5(
        data2[4]), .IN6(n6), .Q(data_o[4]) );
  AO222X1 U10 ( .IN1(data1[3]), .IN2(n8), .IN3(data0[3]), .IN4(n7), .IN5(
        data2[3]), .IN6(n6), .Q(data_o[3]) );
  AO222X1 U11 ( .IN1(data1[2]), .IN2(n8), .IN3(data0[2]), .IN4(n7), .IN5(
        data2[2]), .IN6(n6), .Q(data_o[2]) );
  AO222X1 U12 ( .IN1(data1[1]), .IN2(n8), .IN3(data0[1]), .IN4(n7), .IN5(
        data2[1]), .IN6(n6), .Q(data_o[1]) );
  AO222X1 U13 ( .IN1(data1[15]), .IN2(n8), .IN3(data0[15]), .IN4(n7), .IN5(
        data2[15]), .IN6(n6), .Q(data_o[15]) );
  AO222X1 U14 ( .IN1(data1[14]), .IN2(n8), .IN3(data0[14]), .IN4(n7), .IN5(
        data2[14]), .IN6(n6), .Q(data_o[14]) );
  AO222X1 U15 ( .IN1(data1[13]), .IN2(n8), .IN3(data0[13]), .IN4(n7), .IN5(
        data2[13]), .IN6(n6), .Q(data_o[13]) );
  AO222X1 U16 ( .IN1(data1[12]), .IN2(n8), .IN3(data0[12]), .IN4(n7), .IN5(
        data2[12]), .IN6(n6), .Q(data_o[12]) );
  AO222X1 U17 ( .IN1(data1[11]), .IN2(n8), .IN3(data0[11]), .IN4(n7), .IN5(
        data2[11]), .IN6(n6), .Q(data_o[11]) );
  AO222X1 U18 ( .IN1(data1[10]), .IN2(n8), .IN3(data0[10]), .IN4(n7), .IN5(
        data2[10]), .IN6(n6), .Q(data_o[10]) );
  AO222X1 U19 ( .IN1(data1[0]), .IN2(n8), .IN3(data0[0]), .IN4(n7), .IN5(
        data2[0]), .IN6(n6), .Q(data_o[0]) );
  INVX0 U2 ( .INP(select0), .ZN(n2) );
  INVX0 U3 ( .INP(select1), .ZN(n1) );
  AND3X1 U20 ( .IN1(n2), .IN2(n1), .IN3(select2), .Q(n6) );
  NOR3X0 U21 ( .IN1(select1), .IN2(select2), .IN3(n2), .QN(n7) );
  NOR3X0 U22 ( .IN1(select0), .IN2(select2), .IN3(n1), .QN(n8) );
endmodule



    module node4_NODE_X2_NODE_Y0I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__I_node_2_node_interface__ ( 
        \clk.clk , \reset.reset , \local_node.clk , 
        \local_node.buffer_full_in , \local_node.buffer_full_out , 
        \local_node.receiving_data , \local_node.sending_data , 
        \local_node.data_in , \local_node.data_out , \node_0.clk , 
        \node_0.buffer_full_in , \node_0.buffer_full_out , 
        \node_0.receiving_data , \node_0.sending_data , \node_0.data_in , 
        \node_0.data_out , \node_1.clk , \node_1.buffer_full_in , 
        \node_1.buffer_full_out , \node_1.receiving_data , 
        \node_1.sending_data , \node_1.data_in , \node_1.data_out , 
        \node_2.clk , \node_2.buffer_full_in , \node_2.buffer_full_out , 
        \node_2.receiving_data , \node_2.sending_data , \node_2.data_in , 
        \node_2.data_out  );
  input [15:0] \local_node.data_in ;
  output [15:0] \local_node.data_out ;
  input [15:0] \node_0.data_in ;
  output [15:0] \node_0.data_out ;
  input [15:0] \node_1.data_in ;
  output [15:0] \node_1.data_out ;
  input [15:0] \node_2.data_in ;
  output [15:0] \node_2.data_out ;
  input \clk.clk , \reset.reset , \local_node.buffer_full_in ,
         \local_node.receiving_data , \node_0.buffer_full_in ,
         \node_0.receiving_data , \node_1.buffer_full_in ,
         \node_1.receiving_data , \node_2.buffer_full_in ,
         \node_2.receiving_data ;
  output \local_node.buffer_full_out , \local_node.sending_data ,
         \node_0.buffer_full_out , \node_0.sending_data ,
         \node_1.buffer_full_out , \node_1.sending_data ,
         \node_2.buffer_full_out , \node_2.sending_data ;
  inout \local_node.clk ,  \node_0.clk ,  \node_1.clk ,  \node_2.clk ;
  wire   \buffer_out[3][15] , \buffer_out[3][14] , \buffer_out[3][13] ,
         \buffer_out[3][12] , \buffer_out[3][11] , \buffer_out[3][10] ,
         \buffer_out[3][9] , \buffer_out[3][8] , \buffer_out[3][7] ,
         \buffer_out[3][6] , \buffer_out[3][5] , \buffer_out[3][4] ,
         \buffer_out[3][3] , \buffer_out[3][2] , \buffer_out[3][1] ,
         \buffer_out[3][0] , \buffer_out[2][15] , \buffer_out[2][14] ,
         \buffer_out[2][13] , \buffer_out[2][12] , \buffer_out[2][11] ,
         \buffer_out[2][10] , \buffer_out[2][9] , \buffer_out[2][8] ,
         \buffer_out[2][7] , \buffer_out[2][6] , \buffer_out[2][5] ,
         \buffer_out[2][4] , \buffer_out[2][3] , \buffer_out[2][2] ,
         \buffer_out[2][1] , \buffer_out[2][0] , \buffer_out[1][15] ,
         \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] ,
         \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] ,
         \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] ,
         \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] ,
         \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] ,
         \buffer_out[0][15] , \buffer_out[0][14] , \buffer_out[0][13] ,
         \buffer_out[0][12] , \buffer_out[0][11] , \buffer_out[0][10] ,
         \buffer_out[0][9] , \buffer_out[0][8] , \buffer_out[0][7] ,
         \buffer_out[0][6] , \buffer_out[0][5] , \buffer_out[0][4] ,
         \buffer_out[0][3] , \buffer_out[0][2] , \buffer_out[0][1] ,
         \buffer_out[0][0] , \next_buffer_out[3][15] ,
         \next_buffer_out[3][14] , \next_buffer_out[3][13] ,
         \next_buffer_out[3][12] , \next_buffer_out[3][11] ,
         \next_buffer_out[3][10] , \next_buffer_out[3][9] ,
         \next_buffer_out[3][8] , \next_buffer_out[3][7] ,
         \next_buffer_out[3][6] , \next_buffer_out[3][5] ,
         \next_buffer_out[3][4] , \next_buffer_out[3][3] ,
         \next_buffer_out[3][2] , \next_buffer_out[3][1] ,
         \next_buffer_out[3][0] , \next_buffer_out[2][15] ,
         \next_buffer_out[2][14] , \next_buffer_out[2][13] ,
         \next_buffer_out[2][12] , \next_buffer_out[2][11] ,
         \next_buffer_out[2][10] , \next_buffer_out[2][9] ,
         \next_buffer_out[2][8] , \next_buffer_out[2][7] ,
         \next_buffer_out[2][6] , \next_buffer_out[2][5] ,
         \next_buffer_out[2][4] , \next_buffer_out[2][3] ,
         \next_buffer_out[2][2] , \next_buffer_out[2][1] ,
         \next_buffer_out[2][0] , \next_buffer_out[1][15] ,
         \next_buffer_out[1][14] , \next_buffer_out[1][13] ,
         \next_buffer_out[1][12] , \next_buffer_out[1][11] ,
         \next_buffer_out[1][10] , \next_buffer_out[1][9] ,
         \next_buffer_out[1][8] , \next_buffer_out[1][7] ,
         \next_buffer_out[1][6] , \next_buffer_out[1][5] ,
         \next_buffer_out[1][4] , \next_buffer_out[1][3] ,
         \next_buffer_out[1][2] , \next_buffer_out[1][1] ,
         \next_buffer_out[1][0] , \next_buffer_out[0][15] ,
         \next_buffer_out[0][14] , \next_buffer_out[0][13] ,
         \next_buffer_out[0][12] , \next_buffer_out[0][11] ,
         \next_buffer_out[0][10] , \next_buffer_out[0][9] ,
         \next_buffer_out[0][8] , \next_buffer_out[0][7] ,
         \next_buffer_out[0][6] , \next_buffer_out[0][5] ,
         \next_buffer_out[0][4] , \next_buffer_out[0][3] ,
         \next_buffer_out[0][2] , \next_buffer_out[0][1] ,
         \next_buffer_out[0][0] ;
  wire   [3:0] buffer_full_in;
  wire   [3:0] receiving_data;
  wire   [3:0] pop_v;
  wire   [3:0] data_valid;
  wire   [3:0] next_data_valid;
  wire   [2:0] grant_1;
  wire   [2:0] grant_2;
  wire   [2:0] grant_3;
  tri   \local_node.buffer_full_in ;
  tri   \local_node.buffer_full_out ;
  tri   \local_node.receiving_data ;
  tri   \local_node.sending_data ;
  tri   [15:0] \local_node.data_in ;
  tri   [15:0] \local_node.data_out ;

  converter_out_I_n_node_interface_dut_ c3 ( .\n.buffer_full_in (
        \local_node.buffer_full_in ), .\n.receiving_data (
        \local_node.receiving_data ), .\n.data_in (\local_node.data_in ), 
        .\n.buffer_full_out (\local_node.buffer_full_out ), .\n.sending_data (
        \local_node.sending_data ), .\n.data_out (\local_node.data_out ), 
        .buffer_full_in(1'b0), .receiving_data(1'b0), .data_in({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  fifo_kev_47 \genblk1[0].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[0]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[0]), .data_out({\buffer_out[0][15] , 
        \buffer_out[0][14] , \buffer_out[0][13] , \buffer_out[0][12] , 
        \buffer_out[0][11] , \buffer_out[0][10] , \buffer_out[0][9] , 
        \buffer_out[0][8] , \buffer_out[0][7] , \buffer_out[0][6] , 
        \buffer_out[0][5] , \buffer_out[0][4] , \buffer_out[0][3] , 
        \buffer_out[0][2] , \buffer_out[0][1] , \buffer_out[0][0] }), 
        .next_data_out({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] , 
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .next_data_valid(
        next_data_valid[0]) );
  address_counter_47 \genblk1[0].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] }), 
        .buffer_data_valid(next_data_valid[0]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .buffer_pop(
        pop_v[0]), .receiving_data(1'b0) );
  fifo_kev_46 \genblk1[1].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[1]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[1]), .data_out({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), 
        .next_data_out({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] , 
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .next_data_valid(
        next_data_valid[1]) );
  address_counter_46 \genblk1[1].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] }), 
        .buffer_data_valid(next_data_valid[1]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .buffer_pop(
        pop_v[1]), .receiving_data(1'b0) );
  fifo_kev_45 \genblk1[2].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[2]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[2]), .data_out({\buffer_out[2][15] , 
        \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] , 
        \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] , 
        \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] , 
        \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] , 
        \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] }), 
        .next_data_out({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] , 
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .next_data_valid(
        next_data_valid[2]) );
  address_counter_45 \genblk1[2].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] }), 
        .buffer_data_valid(next_data_valid[2]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .buffer_pop(
        pop_v[2]), .receiving_data(1'b0) );
  fifo_kev_44 \genblk1[3].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[3]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[3]), .data_out({\buffer_out[3][15] , 
        \buffer_out[3][14] , \buffer_out[3][13] , \buffer_out[3][12] , 
        \buffer_out[3][11] , \buffer_out[3][10] , \buffer_out[3][9] , 
        \buffer_out[3][8] , \buffer_out[3][7] , \buffer_out[3][6] , 
        \buffer_out[3][5] , \buffer_out[3][4] , \buffer_out[3][3] , 
        \buffer_out[3][2] , \buffer_out[3][1] , \buffer_out[3][0] }), 
        .next_data_out({\next_buffer_out[3][15] , \next_buffer_out[3][14] , 
        \next_buffer_out[3][13] , \next_buffer_out[3][12] , 
        \next_buffer_out[3][11] , \next_buffer_out[3][10] , 
        \next_buffer_out[3][9] , \next_buffer_out[3][8] , 
        \next_buffer_out[3][7] , \next_buffer_out[3][6] , 
        \next_buffer_out[3][5] , \next_buffer_out[3][4] , 
        \next_buffer_out[3][3] , \next_buffer_out[3][2] , 
        \next_buffer_out[3][1] , \next_buffer_out[3][0] }), .next_data_valid(
        next_data_valid[3]) );
  address_counter_44 \genblk1[3].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[3][15] , \next_buffer_out[3][14] , 
        \next_buffer_out[3][13] , \next_buffer_out[3][12] , 
        \next_buffer_out[3][11] , \next_buffer_out[3][10] , 
        \next_buffer_out[3][9] , \next_buffer_out[3][8] }), 
        .buffer_data_valid(next_data_valid[3]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[3][7] , \next_buffer_out[3][6] , 
        \next_buffer_out[3][5] , \next_buffer_out[3][4] , 
        \next_buffer_out[3][3] , \next_buffer_out[3][2] , 
        \next_buffer_out[3][1] , \next_buffer_out[3][0] }), .buffer_pop(
        pop_v[3]), .receiving_data(1'b0) );
  converter_out_I_n_node_interface_dut_ \genblk2.c0  ( .\n.buffer_full_in (
        \node_0.buffer_full_in ), .\n.receiving_data (\node_0.receiving_data ), 
        .\n.data_in (\node_0.data_in ), .\n.buffer_full_out (
        \node_0.buffer_full_out ), .\n.sending_data (\node_0.sending_data ), 
        .\n.data_out (\node_0.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_in_I_n_node_interface_dut__18 \genblk2.c1  ( .\n.buffer_full_in (
        \node_1.buffer_full_in ), .\n.receiving_data (\node_1.receiving_data ), 
        .\n.data_in (\node_1.data_in ), .\n.buffer_full_out (
        \node_1.buffer_full_out ), .\n.sending_data (\node_1.sending_data ), 
        .\n.data_out (\node_1.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_out_I_n_node_interface_dut_ \genblk2.c2  ( .\n.buffer_full_in (
        \node_2.buffer_full_in ), .\n.receiving_data (\node_2.receiving_data ), 
        .\n.data_in (\node_2.data_in ), .\n.buffer_full_out (
        \node_2.buffer_full_out ), .\n.sending_data (\node_2.sending_data ), 
        .\n.data_out (\node_2.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  controller4_edge_n_0 \genblk2.n  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .packet_addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .local_addr({1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .packet_valid(data_valid), .buffer_full_in({1'b0, 1'b0, 1'b0, 1'b0}), 
        .grant_1(grant_1), .grant_2(grant_2), .grant_3(grant_3), .pop_v(pop_v)
         );
  mux3_1_16 \genblk2.mux_e  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[2][15] , 
        \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] , 
        \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] , 
        \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] , 
        \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] , 
        \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] }), .data2({
        \buffer_out[3][15] , \buffer_out[3][14] , \buffer_out[3][13] , 
        \buffer_out[3][12] , \buffer_out[3][11] , \buffer_out[3][10] , 
        \buffer_out[3][9] , \buffer_out[3][8] , \buffer_out[3][7] , 
        \buffer_out[3][6] , \buffer_out[3][5] , \buffer_out[3][4] , 
        \buffer_out[3][3] , \buffer_out[3][2] , \buffer_out[3][1] , 
        \buffer_out[3][0] }), .select0(grant_1[0]), .select1(grant_1[1]), 
        .select2(grant_1[2]) );
  mux3_1_15 \genblk2.mux_w  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[3][15] , \buffer_out[3][14] , \buffer_out[3][13] , 
        \buffer_out[3][12] , \buffer_out[3][11] , \buffer_out[3][10] , 
        \buffer_out[3][9] , \buffer_out[3][8] , \buffer_out[3][7] , 
        \buffer_out[3][6] , \buffer_out[3][5] , \buffer_out[3][4] , 
        \buffer_out[3][3] , \buffer_out[3][2] , \buffer_out[3][1] , 
        \buffer_out[3][0] }), .select0(grant_2[0]), .select1(grant_2[1]), 
        .select2(grant_2[2]) );
  mux3_1_14 \genblk2.mux_l  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[2][15] , \buffer_out[2][14] , \buffer_out[2][13] , 
        \buffer_out[2][12] , \buffer_out[2][11] , \buffer_out[2][10] , 
        \buffer_out[2][9] , \buffer_out[2][8] , \buffer_out[2][7] , 
        \buffer_out[2][6] , \buffer_out[2][5] , \buffer_out[2][4] , 
        \buffer_out[2][3] , \buffer_out[2][2] , \buffer_out[2][1] , 
        \buffer_out[2][0] }), .select0(grant_3[0]), .select1(grant_3[1]), 
        .select2(grant_3[2]) );
endmodule


module fifo_kev_43 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_87 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_43 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_87 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_86 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_43 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_86 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_43_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_43 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_43 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_43 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_43_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_42 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_85 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_42 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_85 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_84 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_42 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_84 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_42_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_42 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_42 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_42 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_42_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_41 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_83 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_41 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_83 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_82 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_41 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_82 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_41_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_41 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_41 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_41 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_41_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_40 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_81 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_40 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_81 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_80 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_40 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_80 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_40_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_40 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_40 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_40 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_40_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module converter_in_I_n_node_interface_dut__17 ( \n.buffer_full_in , 
        \n.receiving_data , \n.data_in , \n.buffer_full_out , \n.sending_data , 
        \n.data_out , buffer_full_out, sending_data, data_out, buffer_full_in, 
        receiving_data, data_in );
  input [15:0] \n.data_in ;
  output [15:0] \n.data_out ;
  output [15:0] data_out;
  input [15:0] data_in;
  input \n.buffer_full_in , \n.receiving_data , buffer_full_in, receiving_data;
  output \n.buffer_full_out , \n.sending_data , buffer_full_out, sending_data;
  wire   \n.buffer_full_in , \n.receiving_data , buffer_full_in,
         receiving_data;
  assign buffer_full_out = \n.buffer_full_in ;
  assign sending_data = \n.receiving_data ;
  assign data_out[15] = \n.data_in  [15];
  assign data_out[14] = \n.data_in  [14];
  assign data_out[13] = \n.data_in  [13];
  assign data_out[12] = \n.data_in  [12];
  assign data_out[11] = \n.data_in  [11];
  assign data_out[10] = \n.data_in  [10];
  assign data_out[9] = \n.data_in  [9];
  assign data_out[8] = \n.data_in  [8];
  assign data_out[7] = \n.data_in  [7];
  assign data_out[6] = \n.data_in  [6];
  assign data_out[5] = \n.data_in  [5];
  assign data_out[4] = \n.data_in  [4];
  assign data_out[3] = \n.data_in  [3];
  assign data_out[2] = \n.data_in  [2];
  assign data_out[1] = \n.data_in  [1];
  assign data_out[0] = \n.data_in  [0];
  assign \n.buffer_full_out  = buffer_full_in;
  assign \n.sending_data  = receiving_data;
  assign \n.data_out  [15] = data_in[15];
  assign \n.data_out  [14] = data_in[14];
  assign \n.data_out  [13] = data_in[13];
  assign \n.data_out  [12] = data_in[12];
  assign \n.data_out  [11] = data_in[11];
  assign \n.data_out  [10] = data_in[10];
  assign \n.data_out  [9] = data_in[9];
  assign \n.data_out  [8] = data_in[8];
  assign \n.data_out  [7] = data_in[7];
  assign \n.data_out  [6] = data_in[6];
  assign \n.data_out  [5] = data_in[5];
  assign \n.data_out  [4] = data_in[4];
  assign \n.data_out  [3] = data_in[3];
  assign \n.data_out  [2] = data_in[2];
  assign \n.data_out  [1] = data_in[1];
  assign \n.data_out  [0] = data_in[0];

endmodule


module converter_in_I_n_node_interface_dut__16 ( \n.buffer_full_in , 
        \n.receiving_data , \n.data_in , \n.buffer_full_out , \n.sending_data , 
        \n.data_out , buffer_full_out, sending_data, data_out, buffer_full_in, 
        receiving_data, data_in );
  input [15:0] \n.data_in ;
  output [15:0] \n.data_out ;
  output [15:0] data_out;
  input [15:0] data_in;
  input \n.buffer_full_in , \n.receiving_data , buffer_full_in, receiving_data;
  output \n.buffer_full_out , \n.sending_data , buffer_full_out, sending_data;
  wire   \n.buffer_full_in , \n.receiving_data , buffer_full_in,
         receiving_data;
  assign buffer_full_out = \n.buffer_full_in ;
  assign sending_data = \n.receiving_data ;
  assign data_out[15] = \n.data_in  [15];
  assign data_out[14] = \n.data_in  [14];
  assign data_out[13] = \n.data_in  [13];
  assign data_out[12] = \n.data_in  [12];
  assign data_out[11] = \n.data_in  [11];
  assign data_out[10] = \n.data_in  [10];
  assign data_out[9] = \n.data_in  [9];
  assign data_out[8] = \n.data_in  [8];
  assign data_out[7] = \n.data_in  [7];
  assign data_out[6] = \n.data_in  [6];
  assign data_out[5] = \n.data_in  [5];
  assign data_out[4] = \n.data_in  [4];
  assign data_out[3] = \n.data_in  [3];
  assign data_out[2] = \n.data_in  [2];
  assign data_out[1] = \n.data_in  [1];
  assign data_out[0] = \n.data_in  [0];
  assign \n.buffer_full_out  = buffer_full_in;
  assign \n.sending_data  = receiving_data;
  assign \n.data_out  [15] = data_in[15];
  assign \n.data_out  [14] = data_in[14];
  assign \n.data_out  [13] = data_in[13];
  assign \n.data_out  [12] = data_in[12];
  assign \n.data_out  [11] = data_in[11];
  assign \n.data_out  [10] = data_in[10];
  assign \n.data_out  [9] = data_in[9];
  assign \n.data_out  [8] = data_in[8];
  assign \n.data_out  [7] = data_in[7];
  assign \n.data_out  [6] = data_in[6];
  assign \n.data_out  [5] = data_in[5];
  assign \n.data_out  [4] = data_in[4];
  assign \n.data_out  [3] = data_in[3];
  assign \n.data_out  [2] = data_in[2];
  assign \n.data_out  [1] = data_in[1];
  assign \n.data_out  [0] = data_in[0];

endmodule


module flipflop_BITS3_27 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_27 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_27 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS3_26 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_26 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_26 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS1_67 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_67 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_67 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_66 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_66 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_66 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter3_13 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [2:0] request;
  output [2:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[1][2] , \req_i[1][1] , \req_i[1][0] , \req_i[0][2] ,
         \req_i[0][1] , tail_en, N99, N100, N101, N110, N111, N118, N119, N120,
         N121, n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [1:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N99 = request[0];
  assign N100 = request[1];
  assign N101 = request[2];

  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(N111), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(N110), .Q(\req_i[0][1] ) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N121), .D(tail_en), .Q(req_en[0]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N120), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N119), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N118), .Q(grant[0]) );
  AND2X1 U20 ( .IN1(n8), .IN2(N101), .Q(n7) );
  OR3X1 U21 ( .IN1(n3), .IN2(N111), .IN3(n6), .Q(N121) );
  NOR3X0 U22 ( .IN1(N99), .IN2(N100), .IN3(n6), .QN(N120) );
  NOR3X0 U23 ( .IN1(n2), .IN2(N99), .IN3(n6), .QN(N119) );
  NAND3X0 U24 ( .IN1(n2), .IN2(n3), .IN3(n1), .QN(n5) );
  AO22X1 U25 ( .IN1(N100), .IN2(N101), .IN3(N99), .IN4(N101), .Q(N111) );
  INVX0 U10 ( .INP(N101), .ZN(n3) );
  NAND2X1 U11 ( .IN1(n5), .IN2(n4), .QN(n6) );
  INVX0 U12 ( .INP(N99), .ZN(n1) );
  INVX0 U13 ( .INP(N100), .ZN(n2) );
  INVX0 U14 ( .INP(buffer_full_i), .ZN(n4) );
  NAND2X1 U15 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NOR2X0 U16 ( .IN1(n1), .IN2(n6), .QN(N118) );
  NOR2X0 U17 ( .IN1(n1), .IN2(n2), .QN(N110) );
  OA21X1 U18 ( .IN1(N110), .IN2(n7), .IN3(n4), .Q(tail_en) );
  OA21X1 U19 ( .IN1(N101), .IN2(n8), .IN3(n4), .Q(grant_v_o) );
  register_BITS3_27 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][2] , \req_i[0][1] , 1'b0}), .data_o({
        1'b0, 1'b0, 1'b0}) );
  register_BITS3_26 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][2] , \req_i[1][1] , \req_i[1][0] }), 
        .data_o({1'b0, 1'b0, 1'b0}) );
  register_BITS1_67 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b1), .data_o(1'b0) );
  register_BITS1_66 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module flipflop_BITS3_25 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_25 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_25 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS3_24 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_24 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_24 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS1_65 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_65 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_65 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_64 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_64 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_64 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter3_12 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [2:0] request;
  output [2:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[1][2] , \req_i[1][1] , \req_i[1][0] , \req_i[0][2] ,
         \req_i[0][1] , tail_en, N99, N100, N101, N110, N111, N118, N119, N120,
         N121, n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [1:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N99 = request[0];
  assign N100 = request[1];
  assign N101 = request[2];

  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(N111), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(N110), .Q(\req_i[0][1] ) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N121), .D(tail_en), .Q(req_en[0]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N120), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N119), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N118), .Q(grant[0]) );
  AND2X1 U20 ( .IN1(n8), .IN2(N101), .Q(n7) );
  OR3X1 U21 ( .IN1(n3), .IN2(N111), .IN3(n6), .Q(N121) );
  NOR3X0 U22 ( .IN1(N99), .IN2(N100), .IN3(n6), .QN(N120) );
  NOR3X0 U23 ( .IN1(n2), .IN2(N99), .IN3(n6), .QN(N119) );
  NAND3X0 U24 ( .IN1(n2), .IN2(n3), .IN3(n1), .QN(n5) );
  AO22X1 U25 ( .IN1(N100), .IN2(N101), .IN3(N99), .IN4(N101), .Q(N111) );
  INVX0 U10 ( .INP(N101), .ZN(n3) );
  NAND2X1 U11 ( .IN1(n5), .IN2(n4), .QN(n6) );
  INVX0 U12 ( .INP(N99), .ZN(n1) );
  INVX0 U13 ( .INP(N100), .ZN(n2) );
  INVX0 U14 ( .INP(buffer_full_i), .ZN(n4) );
  NAND2X1 U15 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NOR2X0 U16 ( .IN1(n1), .IN2(n6), .QN(N118) );
  NOR2X0 U17 ( .IN1(n1), .IN2(n2), .QN(N110) );
  OA21X1 U18 ( .IN1(N110), .IN2(n7), .IN3(n4), .Q(tail_en) );
  OA21X1 U19 ( .IN1(N101), .IN2(n8), .IN3(n4), .Q(grant_v_o) );
  register_BITS3_25 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][2] , \req_i[0][1] , 1'b0}), .data_o({
        1'b0, 1'b0, 1'b0}) );
  register_BITS3_24 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][2] , \req_i[1][1] , \req_i[1][0] }), 
        .data_o({1'b0, 1'b0, 1'b0}) );
  register_BITS1_65 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b1), .data_o(1'b0) );
  register_BITS1_64 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module flipflop_BITS3_23 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_23 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_23 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS3_22 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_22 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_22 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS1_63 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_63 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_63 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_62 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_62 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_62 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter3_11 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [2:0] request;
  output [2:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[1][2] , \req_i[1][1] , \req_i[1][0] , \req_i[0][2] ,
         \req_i[0][1] , tail_en, N99, N100, N101, N110, N111, N118, N119, N120,
         N121, n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [1:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N99 = request[0];
  assign N100 = request[1];
  assign N101 = request[2];

  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(N111), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(N110), .Q(\req_i[0][1] ) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N121), .D(tail_en), .Q(req_en[0]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N120), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N119), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N118), .Q(grant[0]) );
  AND2X1 U20 ( .IN1(n8), .IN2(N101), .Q(n7) );
  OR3X1 U21 ( .IN1(n3), .IN2(N111), .IN3(n6), .Q(N121) );
  NOR3X0 U22 ( .IN1(N99), .IN2(N100), .IN3(n6), .QN(N120) );
  NOR3X0 U23 ( .IN1(n2), .IN2(N99), .IN3(n6), .QN(N119) );
  NAND3X0 U24 ( .IN1(n2), .IN2(n3), .IN3(n1), .QN(n5) );
  AO22X1 U25 ( .IN1(N100), .IN2(N101), .IN3(N99), .IN4(N101), .Q(N111) );
  INVX0 U10 ( .INP(N101), .ZN(n3) );
  NAND2X1 U11 ( .IN1(n5), .IN2(n4), .QN(n6) );
  INVX0 U12 ( .INP(N99), .ZN(n1) );
  INVX0 U13 ( .INP(N100), .ZN(n2) );
  INVX0 U14 ( .INP(buffer_full_i), .ZN(n4) );
  NAND2X1 U15 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NOR2X0 U16 ( .IN1(n1), .IN2(n6), .QN(N118) );
  NOR2X0 U17 ( .IN1(n1), .IN2(n2), .QN(N110) );
  OA21X1 U18 ( .IN1(N110), .IN2(n7), .IN3(n4), .Q(tail_en) );
  OA21X1 U19 ( .IN1(N101), .IN2(n8), .IN3(n4), .Q(grant_v_o) );
  register_BITS3_23 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][2] , \req_i[0][1] , 1'b0}), .data_o({
        1'b0, 1'b0, 1'b0}) );
  register_BITS3_22 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][2] , \req_i[1][1] , \req_i[1][0] }), 
        .data_o({1'b0, 1'b0, 1'b0}) );
  register_BITS1_63 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b1), .data_o(1'b0) );
  register_BITS1_62 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module dccl_43 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_42 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_41 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_40 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module controller4_edge_s_1 ( clk, rst, .packet_addr({\packet_addr[3][7] , 
        \packet_addr[3][6] , \packet_addr[3][5] , \packet_addr[3][4] , 
        \packet_addr[3][3] , \packet_addr[3][2] , \packet_addr[3][1] , 
        \packet_addr[3][0] , \packet_addr[2][7] , \packet_addr[2][6] , 
        \packet_addr[2][5] , \packet_addr[2][4] , \packet_addr[2][3] , 
        \packet_addr[2][2] , \packet_addr[2][1] , \packet_addr[2][0] , 
        \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] , 
        \packet_addr[1][4] , \packet_addr[1][3] , \packet_addr[1][2] , 
        \packet_addr[1][1] , \packet_addr[1][0] , \packet_addr[0][7] , 
        \packet_addr[0][6] , \packet_addr[0][5] , \packet_addr[0][4] , 
        \packet_addr[0][3] , \packet_addr[0][2] , \packet_addr[0][1] , 
        \packet_addr[0][0] }), local_addr, packet_valid, buffer_full_in, 
        grant_1, grant_2, grant_3, grant_v, pop_v );
  input [7:0] local_addr;
  input [3:0] packet_valid;
  input [3:0] buffer_full_in;
  output [2:0] grant_1;
  output [2:0] grant_2;
  output [2:0] grant_3;
  output [3:0] grant_v;
  output [3:0] pop_v;
  input clk, rst, \packet_addr[3][7] , \packet_addr[3][6] ,
         \packet_addr[3][5] , \packet_addr[3][4] , \packet_addr[3][3] ,
         \packet_addr[3][2] , \packet_addr[3][1] , \packet_addr[3][0] ,
         \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] ,
         \packet_addr[2][4] , \packet_addr[2][3] , \packet_addr[2][2] ,
         \packet_addr[2][1] , \packet_addr[2][0] , \packet_addr[1][7] ,
         \packet_addr[1][6] , \packet_addr[1][5] , \packet_addr[1][4] ,
         \packet_addr[1][3] , \packet_addr[1][2] , \packet_addr[1][1] ,
         \packet_addr[1][0] , \packet_addr[0][7] , \packet_addr[0][6] ,
         \packet_addr[0][5] , \packet_addr[0][4] , \packet_addr[0][3] ,
         \packet_addr[0][2] , \packet_addr[0][1] , \packet_addr[0][0] ;
  wire   \request[3][2] , \request[3][1] , \request[3][0] , \request[2][2] ,
         \request[2][1] , \request[2][0] , \request[1][2] , \request[1][1] ,
         \request[1][0] , \request[0][0] , n1;

  OR3X1 U3 ( .IN1(grant_2[2]), .IN2(grant_1[2]), .IN3(grant_v[0]), .Q(pop_v[3]) );
  OR2X1 U4 ( .IN1(grant_1[1]), .IN2(grant_3[2]), .Q(pop_v[2]) );
  OR2X1 U5 ( .IN1(grant_2[1]), .IN2(grant_3[1]), .Q(pop_v[1]) );
  OR3X1 U6 ( .IN1(grant_3[0]), .IN2(grant_2[0]), .IN3(grant_1[0]), .Q(pop_v[0]) );
  NOR2X0 U1 ( .IN1(n1), .IN2(buffer_full_in[0]), .QN(grant_v[0]) );
  INVX0 U2 ( .INP(\request[0][0] ), .ZN(n1) );
  arbiter3_13 arbiter_e ( .clk(clk), .rst(rst), .request({\request[1][2] , 
        \request[1][1] , \request[1][0] }), .buffer_full_i(buffer_full_in[1]), 
        .grant(grant_1), .grant_v_o(grant_v[1]) );
  arbiter3_12 arbiter_w ( .clk(clk), .rst(rst), .request({\request[2][2] , 
        \request[2][1] , \request[2][0] }), .buffer_full_i(buffer_full_in[2]), 
        .grant(grant_2), .grant_v_o(grant_v[2]) );
  arbiter3_11 arbiter_l ( .clk(clk), .rst(rst), .request({\request[3][2] , 
        \request[3][1] , \request[3][0] }), .buffer_full_i(buffer_full_in[3]), 
        .grant(grant_3), .grant_v_o(grant_v[3]) );
  dccl_43 dccl_n ( .packet_addr_y_i({\packet_addr[0][3] , \packet_addr[0][2] , 
        \packet_addr[0][1] , \packet_addr[0][0] }), .packet_addr_x_i({
        \packet_addr[0][7] , \packet_addr[0][6] , \packet_addr[0][5] , 
        \packet_addr[0][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[0]), 
        .east_req(\request[1][0] ), .west_req(\request[2][0] ), .local_req(
        \request[3][0] ) );
  dccl_42 dccl_e ( .packet_addr_y_i({\packet_addr[1][3] , \packet_addr[1][2] , 
        \packet_addr[1][1] , \packet_addr[1][0] }), .packet_addr_x_i({
        \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] , 
        \packet_addr[1][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[1]), 
        .west_req(\request[2][1] ), .local_req(\request[3][1] ) );
  dccl_41 dccl_w ( .packet_addr_y_i({\packet_addr[2][3] , \packet_addr[2][2] , 
        \packet_addr[2][1] , \packet_addr[2][0] }), .packet_addr_x_i({
        \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] , 
        \packet_addr[2][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[2]), 
        .east_req(\request[1][1] ), .local_req(\request[3][2] ) );
  dccl_40 dccl_l ( .packet_addr_y_i({\packet_addr[3][3] , \packet_addr[3][2] , 
        \packet_addr[3][1] , \packet_addr[3][0] }), .packet_addr_x_i({
        \packet_addr[3][7] , \packet_addr[3][6] , \packet_addr[3][5] , 
        \packet_addr[3][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[3]), 
        .north_req(\request[0][0] ), .east_req(\request[1][2] ), .west_req(
        \request[2][2] ) );
endmodule


module mux3_1_13 ( data0, data1, data2, select0, select1, select2, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  output [15:0] data_o;
  input select0, select1, select2;
  wire   n1, n2, n6, n7, n8;

  AO222X1 U4 ( .IN1(data1[9]), .IN2(n8), .IN3(data0[9]), .IN4(n7), .IN5(
        data2[9]), .IN6(n6), .Q(data_o[9]) );
  AO222X1 U5 ( .IN1(data1[8]), .IN2(n8), .IN3(data0[8]), .IN4(n7), .IN5(
        data2[8]), .IN6(n6), .Q(data_o[8]) );
  AO222X1 U6 ( .IN1(data1[7]), .IN2(n8), .IN3(data0[7]), .IN4(n7), .IN5(
        data2[7]), .IN6(n6), .Q(data_o[7]) );
  AO222X1 U7 ( .IN1(data1[6]), .IN2(n8), .IN3(data0[6]), .IN4(n7), .IN5(
        data2[6]), .IN6(n6), .Q(data_o[6]) );
  AO222X1 U8 ( .IN1(data1[5]), .IN2(n8), .IN3(data0[5]), .IN4(n7), .IN5(
        data2[5]), .IN6(n6), .Q(data_o[5]) );
  AO222X1 U9 ( .IN1(data1[4]), .IN2(n8), .IN3(data0[4]), .IN4(n7), .IN5(
        data2[4]), .IN6(n6), .Q(data_o[4]) );
  AO222X1 U10 ( .IN1(data1[3]), .IN2(n8), .IN3(data0[3]), .IN4(n7), .IN5(
        data2[3]), .IN6(n6), .Q(data_o[3]) );
  AO222X1 U11 ( .IN1(data1[2]), .IN2(n8), .IN3(data0[2]), .IN4(n7), .IN5(
        data2[2]), .IN6(n6), .Q(data_o[2]) );
  AO222X1 U12 ( .IN1(data1[1]), .IN2(n8), .IN3(data0[1]), .IN4(n7), .IN5(
        data2[1]), .IN6(n6), .Q(data_o[1]) );
  AO222X1 U13 ( .IN1(data1[15]), .IN2(n8), .IN3(data0[15]), .IN4(n7), .IN5(
        data2[15]), .IN6(n6), .Q(data_o[15]) );
  AO222X1 U14 ( .IN1(data1[14]), .IN2(n8), .IN3(data0[14]), .IN4(n7), .IN5(
        data2[14]), .IN6(n6), .Q(data_o[14]) );
  AO222X1 U15 ( .IN1(data1[13]), .IN2(n8), .IN3(data0[13]), .IN4(n7), .IN5(
        data2[13]), .IN6(n6), .Q(data_o[13]) );
  AO222X1 U16 ( .IN1(data1[12]), .IN2(n8), .IN3(data0[12]), .IN4(n7), .IN5(
        data2[12]), .IN6(n6), .Q(data_o[12]) );
  AO222X1 U17 ( .IN1(data1[11]), .IN2(n8), .IN3(data0[11]), .IN4(n7), .IN5(
        data2[11]), .IN6(n6), .Q(data_o[11]) );
  AO222X1 U18 ( .IN1(data1[10]), .IN2(n8), .IN3(data0[10]), .IN4(n7), .IN5(
        data2[10]), .IN6(n6), .Q(data_o[10]) );
  AO222X1 U19 ( .IN1(data1[0]), .IN2(n8), .IN3(data0[0]), .IN4(n7), .IN5(
        data2[0]), .IN6(n6), .Q(data_o[0]) );
  INVX0 U2 ( .INP(select0), .ZN(n2) );
  INVX0 U3 ( .INP(select1), .ZN(n1) );
  AND3X1 U20 ( .IN1(n2), .IN2(n1), .IN3(select2), .Q(n6) );
  NOR3X0 U21 ( .IN1(select1), .IN2(select2), .IN3(n2), .QN(n7) );
  NOR3X0 U22 ( .IN1(select0), .IN2(select2), .IN3(n1), .QN(n8) );
endmodule


module mux3_1_12 ( data0, data1, data2, select0, select1, select2, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  output [15:0] data_o;
  input select0, select1, select2;
  wire   n1, n2, n6, n7, n8;

  AO222X1 U4 ( .IN1(data1[9]), .IN2(n8), .IN3(data0[9]), .IN4(n7), .IN5(
        data2[9]), .IN6(n6), .Q(data_o[9]) );
  AO222X1 U5 ( .IN1(data1[8]), .IN2(n8), .IN3(data0[8]), .IN4(n7), .IN5(
        data2[8]), .IN6(n6), .Q(data_o[8]) );
  AO222X1 U6 ( .IN1(data1[7]), .IN2(n8), .IN3(data0[7]), .IN4(n7), .IN5(
        data2[7]), .IN6(n6), .Q(data_o[7]) );
  AO222X1 U7 ( .IN1(data1[6]), .IN2(n8), .IN3(data0[6]), .IN4(n7), .IN5(
        data2[6]), .IN6(n6), .Q(data_o[6]) );
  AO222X1 U8 ( .IN1(data1[5]), .IN2(n8), .IN3(data0[5]), .IN4(n7), .IN5(
        data2[5]), .IN6(n6), .Q(data_o[5]) );
  AO222X1 U9 ( .IN1(data1[4]), .IN2(n8), .IN3(data0[4]), .IN4(n7), .IN5(
        data2[4]), .IN6(n6), .Q(data_o[4]) );
  AO222X1 U10 ( .IN1(data1[3]), .IN2(n8), .IN3(data0[3]), .IN4(n7), .IN5(
        data2[3]), .IN6(n6), .Q(data_o[3]) );
  AO222X1 U11 ( .IN1(data1[2]), .IN2(n8), .IN3(data0[2]), .IN4(n7), .IN5(
        data2[2]), .IN6(n6), .Q(data_o[2]) );
  AO222X1 U12 ( .IN1(data1[1]), .IN2(n8), .IN3(data0[1]), .IN4(n7), .IN5(
        data2[1]), .IN6(n6), .Q(data_o[1]) );
  AO222X1 U13 ( .IN1(data1[15]), .IN2(n8), .IN3(data0[15]), .IN4(n7), .IN5(
        data2[15]), .IN6(n6), .Q(data_o[15]) );
  AO222X1 U14 ( .IN1(data1[14]), .IN2(n8), .IN3(data0[14]), .IN4(n7), .IN5(
        data2[14]), .IN6(n6), .Q(data_o[14]) );
  AO222X1 U15 ( .IN1(data1[13]), .IN2(n8), .IN3(data0[13]), .IN4(n7), .IN5(
        data2[13]), .IN6(n6), .Q(data_o[13]) );
  AO222X1 U16 ( .IN1(data1[12]), .IN2(n8), .IN3(data0[12]), .IN4(n7), .IN5(
        data2[12]), .IN6(n6), .Q(data_o[12]) );
  AO222X1 U17 ( .IN1(data1[11]), .IN2(n8), .IN3(data0[11]), .IN4(n7), .IN5(
        data2[11]), .IN6(n6), .Q(data_o[11]) );
  AO222X1 U18 ( .IN1(data1[10]), .IN2(n8), .IN3(data0[10]), .IN4(n7), .IN5(
        data2[10]), .IN6(n6), .Q(data_o[10]) );
  AO222X1 U19 ( .IN1(data1[0]), .IN2(n8), .IN3(data0[0]), .IN4(n7), .IN5(
        data2[0]), .IN6(n6), .Q(data_o[0]) );
  INVX0 U2 ( .INP(select0), .ZN(n2) );
  INVX0 U3 ( .INP(select1), .ZN(n1) );
  AND3X1 U20 ( .IN1(n2), .IN2(n1), .IN3(select2), .Q(n6) );
  NOR3X0 U21 ( .IN1(select1), .IN2(select2), .IN3(n2), .QN(n7) );
  NOR3X0 U22 ( .IN1(select0), .IN2(select2), .IN3(n1), .QN(n8) );
endmodule


module mux3_1_11 ( data0, data1, data2, select0, select1, select2, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  output [15:0] data_o;
  input select0, select1, select2;
  wire   n1, n2, n6, n7, n8;

  AO222X1 U4 ( .IN1(data1[9]), .IN2(n8), .IN3(data0[9]), .IN4(n7), .IN5(
        data2[9]), .IN6(n6), .Q(data_o[9]) );
  AO222X1 U5 ( .IN1(data1[8]), .IN2(n8), .IN3(data0[8]), .IN4(n7), .IN5(
        data2[8]), .IN6(n6), .Q(data_o[8]) );
  AO222X1 U6 ( .IN1(data1[7]), .IN2(n8), .IN3(data0[7]), .IN4(n7), .IN5(
        data2[7]), .IN6(n6), .Q(data_o[7]) );
  AO222X1 U7 ( .IN1(data1[6]), .IN2(n8), .IN3(data0[6]), .IN4(n7), .IN5(
        data2[6]), .IN6(n6), .Q(data_o[6]) );
  AO222X1 U8 ( .IN1(data1[5]), .IN2(n8), .IN3(data0[5]), .IN4(n7), .IN5(
        data2[5]), .IN6(n6), .Q(data_o[5]) );
  AO222X1 U9 ( .IN1(data1[4]), .IN2(n8), .IN3(data0[4]), .IN4(n7), .IN5(
        data2[4]), .IN6(n6), .Q(data_o[4]) );
  AO222X1 U10 ( .IN1(data1[3]), .IN2(n8), .IN3(data0[3]), .IN4(n7), .IN5(
        data2[3]), .IN6(n6), .Q(data_o[3]) );
  AO222X1 U11 ( .IN1(data1[2]), .IN2(n8), .IN3(data0[2]), .IN4(n7), .IN5(
        data2[2]), .IN6(n6), .Q(data_o[2]) );
  AO222X1 U12 ( .IN1(data1[1]), .IN2(n8), .IN3(data0[1]), .IN4(n7), .IN5(
        data2[1]), .IN6(n6), .Q(data_o[1]) );
  AO222X1 U13 ( .IN1(data1[15]), .IN2(n8), .IN3(data0[15]), .IN4(n7), .IN5(
        data2[15]), .IN6(n6), .Q(data_o[15]) );
  AO222X1 U14 ( .IN1(data1[14]), .IN2(n8), .IN3(data0[14]), .IN4(n7), .IN5(
        data2[14]), .IN6(n6), .Q(data_o[14]) );
  AO222X1 U15 ( .IN1(data1[13]), .IN2(n8), .IN3(data0[13]), .IN4(n7), .IN5(
        data2[13]), .IN6(n6), .Q(data_o[13]) );
  AO222X1 U16 ( .IN1(data1[12]), .IN2(n8), .IN3(data0[12]), .IN4(n7), .IN5(
        data2[12]), .IN6(n6), .Q(data_o[12]) );
  AO222X1 U17 ( .IN1(data1[11]), .IN2(n8), .IN3(data0[11]), .IN4(n7), .IN5(
        data2[11]), .IN6(n6), .Q(data_o[11]) );
  AO222X1 U18 ( .IN1(data1[10]), .IN2(n8), .IN3(data0[10]), .IN4(n7), .IN5(
        data2[10]), .IN6(n6), .Q(data_o[10]) );
  AO222X1 U19 ( .IN1(data1[0]), .IN2(n8), .IN3(data0[0]), .IN4(n7), .IN5(
        data2[0]), .IN6(n6), .Q(data_o[0]) );
  INVX0 U2 ( .INP(select0), .ZN(n2) );
  INVX0 U3 ( .INP(select1), .ZN(n1) );
  AND3X1 U20 ( .IN1(n2), .IN2(n1), .IN3(select2), .Q(n6) );
  NOR3X0 U21 ( .IN1(select1), .IN2(select2), .IN3(n2), .QN(n7) );
  NOR3X0 U22 ( .IN1(select0), .IN2(select2), .IN3(n1), .QN(n8) );
endmodule



    module node4_NODE_X1_NODE_Y3I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__I_node_2_node_interface__ ( 
        \clk.clk , \reset.reset , \local_node.clk , 
        \local_node.buffer_full_in , \local_node.buffer_full_out , 
        \local_node.receiving_data , \local_node.sending_data , 
        \local_node.data_in , \local_node.data_out , \node_0.clk , 
        \node_0.buffer_full_in , \node_0.buffer_full_out , 
        \node_0.receiving_data , \node_0.sending_data , \node_0.data_in , 
        \node_0.data_out , \node_1.clk , \node_1.buffer_full_in , 
        \node_1.buffer_full_out , \node_1.receiving_data , 
        \node_1.sending_data , \node_1.data_in , \node_1.data_out , 
        \node_2.clk , \node_2.buffer_full_in , \node_2.buffer_full_out , 
        \node_2.receiving_data , \node_2.sending_data , \node_2.data_in , 
        \node_2.data_out  );
  input [15:0] \local_node.data_in ;
  output [15:0] \local_node.data_out ;
  input [15:0] \node_0.data_in ;
  output [15:0] \node_0.data_out ;
  input [15:0] \node_1.data_in ;
  output [15:0] \node_1.data_out ;
  input [15:0] \node_2.data_in ;
  output [15:0] \node_2.data_out ;
  input \clk.clk , \reset.reset , \local_node.buffer_full_in ,
         \local_node.receiving_data , \node_0.buffer_full_in ,
         \node_0.receiving_data , \node_1.buffer_full_in ,
         \node_1.receiving_data , \node_2.buffer_full_in ,
         \node_2.receiving_data ;
  output \local_node.buffer_full_out , \local_node.sending_data ,
         \node_0.buffer_full_out , \node_0.sending_data ,
         \node_1.buffer_full_out , \node_1.sending_data ,
         \node_2.buffer_full_out , \node_2.sending_data ;
  inout \local_node.clk ,  \node_0.clk ,  \node_1.clk ,  \node_2.clk ;
  wire   \buffer_out[3][15] , \buffer_out[3][14] , \buffer_out[3][13] ,
         \buffer_out[3][12] , \buffer_out[3][11] , \buffer_out[3][10] ,
         \buffer_out[3][9] , \buffer_out[3][8] , \buffer_out[3][7] ,
         \buffer_out[3][6] , \buffer_out[3][5] , \buffer_out[3][4] ,
         \buffer_out[3][3] , \buffer_out[3][2] , \buffer_out[3][1] ,
         \buffer_out[3][0] , \buffer_out[2][15] , \buffer_out[2][14] ,
         \buffer_out[2][13] , \buffer_out[2][12] , \buffer_out[2][11] ,
         \buffer_out[2][10] , \buffer_out[2][9] , \buffer_out[2][8] ,
         \buffer_out[2][7] , \buffer_out[2][6] , \buffer_out[2][5] ,
         \buffer_out[2][4] , \buffer_out[2][3] , \buffer_out[2][2] ,
         \buffer_out[2][1] , \buffer_out[2][0] , \buffer_out[1][15] ,
         \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] ,
         \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] ,
         \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] ,
         \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] ,
         \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] ,
         \buffer_out[0][15] , \buffer_out[0][14] , \buffer_out[0][13] ,
         \buffer_out[0][12] , \buffer_out[0][11] , \buffer_out[0][10] ,
         \buffer_out[0][9] , \buffer_out[0][8] , \buffer_out[0][7] ,
         \buffer_out[0][6] , \buffer_out[0][5] , \buffer_out[0][4] ,
         \buffer_out[0][3] , \buffer_out[0][2] , \buffer_out[0][1] ,
         \buffer_out[0][0] , \next_buffer_out[3][15] ,
         \next_buffer_out[3][14] , \next_buffer_out[3][13] ,
         \next_buffer_out[3][12] , \next_buffer_out[3][11] ,
         \next_buffer_out[3][10] , \next_buffer_out[3][9] ,
         \next_buffer_out[3][8] , \next_buffer_out[3][7] ,
         \next_buffer_out[3][6] , \next_buffer_out[3][5] ,
         \next_buffer_out[3][4] , \next_buffer_out[3][3] ,
         \next_buffer_out[3][2] , \next_buffer_out[3][1] ,
         \next_buffer_out[3][0] , \next_buffer_out[2][15] ,
         \next_buffer_out[2][14] , \next_buffer_out[2][13] ,
         \next_buffer_out[2][12] , \next_buffer_out[2][11] ,
         \next_buffer_out[2][10] , \next_buffer_out[2][9] ,
         \next_buffer_out[2][8] , \next_buffer_out[2][7] ,
         \next_buffer_out[2][6] , \next_buffer_out[2][5] ,
         \next_buffer_out[2][4] , \next_buffer_out[2][3] ,
         \next_buffer_out[2][2] , \next_buffer_out[2][1] ,
         \next_buffer_out[2][0] , \next_buffer_out[1][15] ,
         \next_buffer_out[1][14] , \next_buffer_out[1][13] ,
         \next_buffer_out[1][12] , \next_buffer_out[1][11] ,
         \next_buffer_out[1][10] , \next_buffer_out[1][9] ,
         \next_buffer_out[1][8] , \next_buffer_out[1][7] ,
         \next_buffer_out[1][6] , \next_buffer_out[1][5] ,
         \next_buffer_out[1][4] , \next_buffer_out[1][3] ,
         \next_buffer_out[1][2] , \next_buffer_out[1][1] ,
         \next_buffer_out[1][0] , \next_buffer_out[0][15] ,
         \next_buffer_out[0][14] , \next_buffer_out[0][13] ,
         \next_buffer_out[0][12] , \next_buffer_out[0][11] ,
         \next_buffer_out[0][10] , \next_buffer_out[0][9] ,
         \next_buffer_out[0][8] , \next_buffer_out[0][7] ,
         \next_buffer_out[0][6] , \next_buffer_out[0][5] ,
         \next_buffer_out[0][4] , \next_buffer_out[0][3] ,
         \next_buffer_out[0][2] , \next_buffer_out[0][1] ,
         \next_buffer_out[0][0] ;
  wire   [3:0] buffer_full_in;
  wire   [3:0] receiving_data;
  wire   [3:0] pop_v;
  wire   [3:0] data_valid;
  wire   [3:0] next_data_valid;
  wire   [2:0] grant_1;
  wire   [2:0] grant_2;
  wire   [2:0] grant_3;
  tri   \local_node.buffer_full_in ;
  tri   \local_node.buffer_full_out ;
  tri   \local_node.receiving_data ;
  tri   \local_node.sending_data ;
  tri   [15:0] \local_node.data_in ;
  tri   [15:0] \local_node.data_out ;

  converter_out_I_n_node_interface_dut_ c3 ( .\n.buffer_full_in (
        \local_node.buffer_full_in ), .\n.receiving_data (
        \local_node.receiving_data ), .\n.data_in (\local_node.data_in ), 
        .\n.buffer_full_out (\local_node.buffer_full_out ), .\n.sending_data (
        \local_node.sending_data ), .\n.data_out (\local_node.data_out ), 
        .buffer_full_in(1'b0), .receiving_data(1'b0), .data_in({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  fifo_kev_43 \genblk1[0].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[0]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[0]), .data_out({\buffer_out[0][15] , 
        \buffer_out[0][14] , \buffer_out[0][13] , \buffer_out[0][12] , 
        \buffer_out[0][11] , \buffer_out[0][10] , \buffer_out[0][9] , 
        \buffer_out[0][8] , \buffer_out[0][7] , \buffer_out[0][6] , 
        \buffer_out[0][5] , \buffer_out[0][4] , \buffer_out[0][3] , 
        \buffer_out[0][2] , \buffer_out[0][1] , \buffer_out[0][0] }), 
        .next_data_out({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] , 
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .next_data_valid(
        next_data_valid[0]) );
  address_counter_43 \genblk1[0].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] }), 
        .buffer_data_valid(next_data_valid[0]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .buffer_pop(
        pop_v[0]), .receiving_data(1'b0) );
  fifo_kev_42 \genblk1[1].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[1]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[1]), .data_out({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), 
        .next_data_out({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] , 
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .next_data_valid(
        next_data_valid[1]) );
  address_counter_42 \genblk1[1].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] }), 
        .buffer_data_valid(next_data_valid[1]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .buffer_pop(
        pop_v[1]), .receiving_data(1'b0) );
  fifo_kev_41 \genblk1[2].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[2]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[2]), .data_out({\buffer_out[2][15] , 
        \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] , 
        \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] , 
        \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] , 
        \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] , 
        \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] }), 
        .next_data_out({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] , 
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .next_data_valid(
        next_data_valid[2]) );
  address_counter_41 \genblk1[2].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] }), 
        .buffer_data_valid(next_data_valid[2]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .buffer_pop(
        pop_v[2]), .receiving_data(1'b0) );
  fifo_kev_40 \genblk1[3].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[3]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[3]), .data_out({\buffer_out[3][15] , 
        \buffer_out[3][14] , \buffer_out[3][13] , \buffer_out[3][12] , 
        \buffer_out[3][11] , \buffer_out[3][10] , \buffer_out[3][9] , 
        \buffer_out[3][8] , \buffer_out[3][7] , \buffer_out[3][6] , 
        \buffer_out[3][5] , \buffer_out[3][4] , \buffer_out[3][3] , 
        \buffer_out[3][2] , \buffer_out[3][1] , \buffer_out[3][0] }), 
        .next_data_out({\next_buffer_out[3][15] , \next_buffer_out[3][14] , 
        \next_buffer_out[3][13] , \next_buffer_out[3][12] , 
        \next_buffer_out[3][11] , \next_buffer_out[3][10] , 
        \next_buffer_out[3][9] , \next_buffer_out[3][8] , 
        \next_buffer_out[3][7] , \next_buffer_out[3][6] , 
        \next_buffer_out[3][5] , \next_buffer_out[3][4] , 
        \next_buffer_out[3][3] , \next_buffer_out[3][2] , 
        \next_buffer_out[3][1] , \next_buffer_out[3][0] }), .next_data_valid(
        next_data_valid[3]) );
  address_counter_40 \genblk1[3].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[3][15] , \next_buffer_out[3][14] , 
        \next_buffer_out[3][13] , \next_buffer_out[3][12] , 
        \next_buffer_out[3][11] , \next_buffer_out[3][10] , 
        \next_buffer_out[3][9] , \next_buffer_out[3][8] }), 
        .buffer_data_valid(next_data_valid[3]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[3][7] , \next_buffer_out[3][6] , 
        \next_buffer_out[3][5] , \next_buffer_out[3][4] , 
        \next_buffer_out[3][3] , \next_buffer_out[3][2] , 
        \next_buffer_out[3][1] , \next_buffer_out[3][0] }), .buffer_pop(
        pop_v[3]), .receiving_data(1'b0) );
  converter_in_I_n_node_interface_dut__17 \genblk2.c0  ( .\n.buffer_full_in (
        \node_0.buffer_full_in ), .\n.receiving_data (\node_0.receiving_data ), 
        .\n.data_in (\node_0.data_in ), .\n.buffer_full_out (
        \node_0.buffer_full_out ), .\n.sending_data (\node_0.sending_data ), 
        .\n.data_out (\node_0.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_in_I_n_node_interface_dut__16 \genblk2.c1  ( .\n.buffer_full_in (
        \node_1.buffer_full_in ), .\n.receiving_data (\node_1.receiving_data ), 
        .\n.data_in (\node_1.data_in ), .\n.buffer_full_out (
        \node_1.buffer_full_out ), .\n.sending_data (\node_1.sending_data ), 
        .\n.data_out (\node_1.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_out_I_n_node_interface_dut_ \genblk2.c2  ( .\n.buffer_full_in (
        \node_2.buffer_full_in ), .\n.receiving_data (\node_2.receiving_data ), 
        .\n.data_in (\node_2.data_in ), .\n.buffer_full_out (
        \node_2.buffer_full_out ), .\n.sending_data (\node_2.sending_data ), 
        .\n.data_out (\node_2.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  controller4_edge_s_1 \genblk2.s  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .packet_addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .local_addr({1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1}), 
        .packet_valid(data_valid), .buffer_full_in({1'b0, 1'b0, 1'b0, 1'b0}), 
        .grant_1(grant_1), .grant_2(grant_2), .grant_3(grant_3), .pop_v(pop_v)
         );
  mux3_1_13 \genblk2.mux_e  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[2][15] , 
        \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] , 
        \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] , 
        \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] , 
        \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] , 
        \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] }), .data2({
        \buffer_out[3][15] , \buffer_out[3][14] , \buffer_out[3][13] , 
        \buffer_out[3][12] , \buffer_out[3][11] , \buffer_out[3][10] , 
        \buffer_out[3][9] , \buffer_out[3][8] , \buffer_out[3][7] , 
        \buffer_out[3][6] , \buffer_out[3][5] , \buffer_out[3][4] , 
        \buffer_out[3][3] , \buffer_out[3][2] , \buffer_out[3][1] , 
        \buffer_out[3][0] }), .select0(grant_1[0]), .select1(grant_1[1]), 
        .select2(grant_1[2]) );
  mux3_1_12 \genblk2.mux_w  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[3][15] , \buffer_out[3][14] , \buffer_out[3][13] , 
        \buffer_out[3][12] , \buffer_out[3][11] , \buffer_out[3][10] , 
        \buffer_out[3][9] , \buffer_out[3][8] , \buffer_out[3][7] , 
        \buffer_out[3][6] , \buffer_out[3][5] , \buffer_out[3][4] , 
        \buffer_out[3][3] , \buffer_out[3][2] , \buffer_out[3][1] , 
        \buffer_out[3][0] }), .select0(grant_2[0]), .select1(grant_2[1]), 
        .select2(grant_2[2]) );
  mux3_1_11 \genblk2.mux_l  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[2][15] , \buffer_out[2][14] , \buffer_out[2][13] , 
        \buffer_out[2][12] , \buffer_out[2][11] , \buffer_out[2][10] , 
        \buffer_out[2][9] , \buffer_out[2][8] , \buffer_out[2][7] , 
        \buffer_out[2][6] , \buffer_out[2][5] , \buffer_out[2][4] , 
        \buffer_out[2][3] , \buffer_out[2][2] , \buffer_out[2][1] , 
        \buffer_out[2][0] }), .select0(grant_3[0]), .select1(grant_3[1]), 
        .select2(grant_3[2]) );
endmodule


module fifo_kev_39 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_79 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_39 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_79 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_78 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_39 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_78 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_39_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_39 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_39 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_39 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_39_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_38 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_77 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_38 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_77 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_76 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_38 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_76 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_38_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_38 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_38 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_38 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_38_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_37 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_75 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_37 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_75 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_74 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_37 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_74 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_37_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_37 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_37 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_37 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_37_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_36 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_73 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_36 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_73 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_72 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_36 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_72 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_36_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_36 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_36 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_36 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_36_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module converter_in_I_n_node_interface_dut__15 ( \n.buffer_full_in , 
        \n.receiving_data , \n.data_in , \n.buffer_full_out , \n.sending_data , 
        \n.data_out , buffer_full_out, sending_data, data_out, buffer_full_in, 
        receiving_data, data_in );
  input [15:0] \n.data_in ;
  output [15:0] \n.data_out ;
  output [15:0] data_out;
  input [15:0] data_in;
  input \n.buffer_full_in , \n.receiving_data , buffer_full_in, receiving_data;
  output \n.buffer_full_out , \n.sending_data , buffer_full_out, sending_data;
  wire   \n.buffer_full_in , \n.receiving_data , buffer_full_in,
         receiving_data;
  assign buffer_full_out = \n.buffer_full_in ;
  assign sending_data = \n.receiving_data ;
  assign data_out[15] = \n.data_in  [15];
  assign data_out[14] = \n.data_in  [14];
  assign data_out[13] = \n.data_in  [13];
  assign data_out[12] = \n.data_in  [12];
  assign data_out[11] = \n.data_in  [11];
  assign data_out[10] = \n.data_in  [10];
  assign data_out[9] = \n.data_in  [9];
  assign data_out[8] = \n.data_in  [8];
  assign data_out[7] = \n.data_in  [7];
  assign data_out[6] = \n.data_in  [6];
  assign data_out[5] = \n.data_in  [5];
  assign data_out[4] = \n.data_in  [4];
  assign data_out[3] = \n.data_in  [3];
  assign data_out[2] = \n.data_in  [2];
  assign data_out[1] = \n.data_in  [1];
  assign data_out[0] = \n.data_in  [0];
  assign \n.buffer_full_out  = buffer_full_in;
  assign \n.sending_data  = receiving_data;
  assign \n.data_out  [15] = data_in[15];
  assign \n.data_out  [14] = data_in[14];
  assign \n.data_out  [13] = data_in[13];
  assign \n.data_out  [12] = data_in[12];
  assign \n.data_out  [11] = data_in[11];
  assign \n.data_out  [10] = data_in[10];
  assign \n.data_out  [9] = data_in[9];
  assign \n.data_out  [8] = data_in[8];
  assign \n.data_out  [7] = data_in[7];
  assign \n.data_out  [6] = data_in[6];
  assign \n.data_out  [5] = data_in[5];
  assign \n.data_out  [4] = data_in[4];
  assign \n.data_out  [3] = data_in[3];
  assign \n.data_out  [2] = data_in[2];
  assign \n.data_out  [1] = data_in[1];
  assign \n.data_out  [0] = data_in[0];

endmodule


module converter_in_I_n_node_interface_dut__14 ( \n.buffer_full_in , 
        \n.receiving_data , \n.data_in , \n.buffer_full_out , \n.sending_data , 
        \n.data_out , buffer_full_out, sending_data, data_out, buffer_full_in, 
        receiving_data, data_in );
  input [15:0] \n.data_in ;
  output [15:0] \n.data_out ;
  output [15:0] data_out;
  input [15:0] data_in;
  input \n.buffer_full_in , \n.receiving_data , buffer_full_in, receiving_data;
  output \n.buffer_full_out , \n.sending_data , buffer_full_out, sending_data;
  wire   \n.buffer_full_in , \n.receiving_data , buffer_full_in,
         receiving_data;
  assign buffer_full_out = \n.buffer_full_in ;
  assign sending_data = \n.receiving_data ;
  assign data_out[15] = \n.data_in  [15];
  assign data_out[14] = \n.data_in  [14];
  assign data_out[13] = \n.data_in  [13];
  assign data_out[12] = \n.data_in  [12];
  assign data_out[11] = \n.data_in  [11];
  assign data_out[10] = \n.data_in  [10];
  assign data_out[9] = \n.data_in  [9];
  assign data_out[8] = \n.data_in  [8];
  assign data_out[7] = \n.data_in  [7];
  assign data_out[6] = \n.data_in  [6];
  assign data_out[5] = \n.data_in  [5];
  assign data_out[4] = \n.data_in  [4];
  assign data_out[3] = \n.data_in  [3];
  assign data_out[2] = \n.data_in  [2];
  assign data_out[1] = \n.data_in  [1];
  assign data_out[0] = \n.data_in  [0];
  assign \n.buffer_full_out  = buffer_full_in;
  assign \n.sending_data  = receiving_data;
  assign \n.data_out  [15] = data_in[15];
  assign \n.data_out  [14] = data_in[14];
  assign \n.data_out  [13] = data_in[13];
  assign \n.data_out  [12] = data_in[12];
  assign \n.data_out  [11] = data_in[11];
  assign \n.data_out  [10] = data_in[10];
  assign \n.data_out  [9] = data_in[9];
  assign \n.data_out  [8] = data_in[8];
  assign \n.data_out  [7] = data_in[7];
  assign \n.data_out  [6] = data_in[6];
  assign \n.data_out  [5] = data_in[5];
  assign \n.data_out  [4] = data_in[4];
  assign \n.data_out  [3] = data_in[3];
  assign \n.data_out  [2] = data_in[2];
  assign \n.data_out  [1] = data_in[1];
  assign \n.data_out  [0] = data_in[0];

endmodule


module flipflop_BITS3_21 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_21 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_21 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS3_20 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_20 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_20 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS1_61 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_61 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_61 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_60 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_60 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_60 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter3_10 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [2:0] request;
  output [2:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[1][2] , \req_i[1][1] , \req_i[1][0] , \req_i[0][2] ,
         \req_i[0][1] , tail_en, N99, N100, N101, N110, N111, N118, N119, N120,
         N121, n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [1:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N99 = request[0];
  assign N100 = request[1];
  assign N101 = request[2];

  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(N111), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(N110), .Q(\req_i[0][1] ) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N121), .D(tail_en), .Q(req_en[0]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N120), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N119), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N118), .Q(grant[0]) );
  AND2X1 U20 ( .IN1(n8), .IN2(N101), .Q(n7) );
  OR3X1 U21 ( .IN1(n3), .IN2(N111), .IN3(n6), .Q(N121) );
  NOR3X0 U22 ( .IN1(N99), .IN2(N100), .IN3(n6), .QN(N120) );
  NOR3X0 U23 ( .IN1(n2), .IN2(N99), .IN3(n6), .QN(N119) );
  NAND3X0 U24 ( .IN1(n2), .IN2(n3), .IN3(n1), .QN(n5) );
  AO22X1 U25 ( .IN1(N100), .IN2(N101), .IN3(N99), .IN4(N101), .Q(N111) );
  INVX0 U10 ( .INP(N101), .ZN(n3) );
  NAND2X1 U11 ( .IN1(n5), .IN2(n4), .QN(n6) );
  INVX0 U12 ( .INP(N99), .ZN(n1) );
  INVX0 U13 ( .INP(N100), .ZN(n2) );
  INVX0 U14 ( .INP(buffer_full_i), .ZN(n4) );
  NAND2X1 U15 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NOR2X0 U16 ( .IN1(n1), .IN2(n6), .QN(N118) );
  NOR2X0 U17 ( .IN1(n1), .IN2(n2), .QN(N110) );
  OA21X1 U18 ( .IN1(N110), .IN2(n7), .IN3(n4), .Q(tail_en) );
  OA21X1 U19 ( .IN1(N101), .IN2(n8), .IN3(n4), .Q(grant_v_o) );
  register_BITS3_21 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][2] , \req_i[0][1] , 1'b0}), .data_o({
        1'b0, 1'b0, 1'b0}) );
  register_BITS3_20 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][2] , \req_i[1][1] , \req_i[1][0] }), 
        .data_o({1'b0, 1'b0, 1'b0}) );
  register_BITS1_61 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b1), .data_o(1'b0) );
  register_BITS1_60 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module flipflop_BITS3_19 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_19 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_19 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS3_18 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_18 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_18 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS1_59 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_59 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_59 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_58 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_58 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_58 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter3_9 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [2:0] request;
  output [2:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[1][2] , \req_i[1][1] , \req_i[1][0] , \req_i[0][2] ,
         \req_i[0][1] , tail_en, N99, N100, N101, N110, N111, N118, N119, N120,
         N121, n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [1:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N99 = request[0];
  assign N100 = request[1];
  assign N101 = request[2];

  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(N111), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(N110), .Q(\req_i[0][1] ) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N121), .D(tail_en), .Q(req_en[0]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N120), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N119), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N118), .Q(grant[0]) );
  AND2X1 U20 ( .IN1(n8), .IN2(N101), .Q(n7) );
  OR3X1 U21 ( .IN1(n3), .IN2(N111), .IN3(n6), .Q(N121) );
  NOR3X0 U22 ( .IN1(N99), .IN2(N100), .IN3(n6), .QN(N120) );
  NOR3X0 U23 ( .IN1(n2), .IN2(N99), .IN3(n6), .QN(N119) );
  NAND3X0 U24 ( .IN1(n2), .IN2(n3), .IN3(n1), .QN(n5) );
  AO22X1 U25 ( .IN1(N100), .IN2(N101), .IN3(N99), .IN4(N101), .Q(N111) );
  INVX0 U10 ( .INP(N101), .ZN(n3) );
  NAND2X1 U11 ( .IN1(n5), .IN2(n4), .QN(n6) );
  INVX0 U12 ( .INP(N99), .ZN(n1) );
  INVX0 U13 ( .INP(N100), .ZN(n2) );
  INVX0 U14 ( .INP(buffer_full_i), .ZN(n4) );
  NAND2X1 U15 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NOR2X0 U16 ( .IN1(n1), .IN2(n6), .QN(N118) );
  NOR2X0 U17 ( .IN1(n1), .IN2(n2), .QN(N110) );
  OA21X1 U18 ( .IN1(N110), .IN2(n7), .IN3(n4), .Q(tail_en) );
  OA21X1 U19 ( .IN1(N101), .IN2(n8), .IN3(n4), .Q(grant_v_o) );
  register_BITS3_19 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][2] , \req_i[0][1] , 1'b0}), .data_o({
        1'b0, 1'b0, 1'b0}) );
  register_BITS3_18 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][2] , \req_i[1][1] , \req_i[1][0] }), 
        .data_o({1'b0, 1'b0, 1'b0}) );
  register_BITS1_59 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b1), .data_o(1'b0) );
  register_BITS1_58 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module flipflop_BITS3_17 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_17 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_17 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS3_16 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_16 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_16 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS1_57 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_57 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_57 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_56 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_56 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_56 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter3_8 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [2:0] request;
  output [2:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[1][2] , \req_i[1][1] , \req_i[1][0] , \req_i[0][2] ,
         \req_i[0][1] , tail_en, N99, N100, N101, N110, N111, N118, N119, N120,
         N121, n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [1:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N99 = request[0];
  assign N100 = request[1];
  assign N101 = request[2];

  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(N111), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(N110), .Q(\req_i[0][1] ) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N121), .D(tail_en), .Q(req_en[0]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N120), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N119), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N118), .Q(grant[0]) );
  AND2X1 U20 ( .IN1(n8), .IN2(N101), .Q(n7) );
  OR3X1 U21 ( .IN1(n3), .IN2(N111), .IN3(n6), .Q(N121) );
  NOR3X0 U22 ( .IN1(N99), .IN2(N100), .IN3(n6), .QN(N120) );
  NOR3X0 U23 ( .IN1(n2), .IN2(N99), .IN3(n6), .QN(N119) );
  NAND3X0 U24 ( .IN1(n2), .IN2(n3), .IN3(n1), .QN(n5) );
  AO22X1 U25 ( .IN1(N100), .IN2(N101), .IN3(N99), .IN4(N101), .Q(N111) );
  INVX0 U10 ( .INP(N101), .ZN(n3) );
  NAND2X1 U11 ( .IN1(n5), .IN2(n4), .QN(n6) );
  INVX0 U12 ( .INP(N99), .ZN(n1) );
  INVX0 U13 ( .INP(N100), .ZN(n2) );
  INVX0 U14 ( .INP(buffer_full_i), .ZN(n4) );
  NAND2X1 U15 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NOR2X0 U16 ( .IN1(n1), .IN2(n6), .QN(N118) );
  NOR2X0 U17 ( .IN1(n1), .IN2(n2), .QN(N110) );
  OA21X1 U18 ( .IN1(N110), .IN2(n7), .IN3(n4), .Q(tail_en) );
  OA21X1 U19 ( .IN1(N101), .IN2(n8), .IN3(n4), .Q(grant_v_o) );
  register_BITS3_17 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][2] , \req_i[0][1] , 1'b0}), .data_o({
        1'b0, 1'b0, 1'b0}) );
  register_BITS3_16 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][2] , \req_i[1][1] , \req_i[1][0] }), 
        .data_o({1'b0, 1'b0, 1'b0}) );
  register_BITS1_57 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b1), .data_o(1'b0) );
  register_BITS1_56 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module dccl_39 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_38 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_37 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_36 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module controller4_edge_s_0 ( clk, rst, .packet_addr({\packet_addr[3][7] , 
        \packet_addr[3][6] , \packet_addr[3][5] , \packet_addr[3][4] , 
        \packet_addr[3][3] , \packet_addr[3][2] , \packet_addr[3][1] , 
        \packet_addr[3][0] , \packet_addr[2][7] , \packet_addr[2][6] , 
        \packet_addr[2][5] , \packet_addr[2][4] , \packet_addr[2][3] , 
        \packet_addr[2][2] , \packet_addr[2][1] , \packet_addr[2][0] , 
        \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] , 
        \packet_addr[1][4] , \packet_addr[1][3] , \packet_addr[1][2] , 
        \packet_addr[1][1] , \packet_addr[1][0] , \packet_addr[0][7] , 
        \packet_addr[0][6] , \packet_addr[0][5] , \packet_addr[0][4] , 
        \packet_addr[0][3] , \packet_addr[0][2] , \packet_addr[0][1] , 
        \packet_addr[0][0] }), local_addr, packet_valid, buffer_full_in, 
        grant_1, grant_2, grant_3, grant_v, pop_v );
  input [7:0] local_addr;
  input [3:0] packet_valid;
  input [3:0] buffer_full_in;
  output [2:0] grant_1;
  output [2:0] grant_2;
  output [2:0] grant_3;
  output [3:0] grant_v;
  output [3:0] pop_v;
  input clk, rst, \packet_addr[3][7] , \packet_addr[3][6] ,
         \packet_addr[3][5] , \packet_addr[3][4] , \packet_addr[3][3] ,
         \packet_addr[3][2] , \packet_addr[3][1] , \packet_addr[3][0] ,
         \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] ,
         \packet_addr[2][4] , \packet_addr[2][3] , \packet_addr[2][2] ,
         \packet_addr[2][1] , \packet_addr[2][0] , \packet_addr[1][7] ,
         \packet_addr[1][6] , \packet_addr[1][5] , \packet_addr[1][4] ,
         \packet_addr[1][3] , \packet_addr[1][2] , \packet_addr[1][1] ,
         \packet_addr[1][0] , \packet_addr[0][7] , \packet_addr[0][6] ,
         \packet_addr[0][5] , \packet_addr[0][4] , \packet_addr[0][3] ,
         \packet_addr[0][2] , \packet_addr[0][1] , \packet_addr[0][0] ;
  wire   \request[3][2] , \request[3][1] , \request[3][0] , \request[2][2] ,
         \request[2][1] , \request[2][0] , \request[1][2] , \request[1][1] ,
         \request[1][0] , \request[0][0] , n1;

  OR3X1 U3 ( .IN1(grant_2[2]), .IN2(grant_1[2]), .IN3(grant_v[0]), .Q(pop_v[3]) );
  OR2X1 U4 ( .IN1(grant_1[1]), .IN2(grant_3[2]), .Q(pop_v[2]) );
  OR2X1 U5 ( .IN1(grant_2[1]), .IN2(grant_3[1]), .Q(pop_v[1]) );
  OR3X1 U6 ( .IN1(grant_3[0]), .IN2(grant_2[0]), .IN3(grant_1[0]), .Q(pop_v[0]) );
  NOR2X0 U1 ( .IN1(n1), .IN2(buffer_full_in[0]), .QN(grant_v[0]) );
  INVX0 U2 ( .INP(\request[0][0] ), .ZN(n1) );
  arbiter3_10 arbiter_e ( .clk(clk), .rst(rst), .request({\request[1][2] , 
        \request[1][1] , \request[1][0] }), .buffer_full_i(buffer_full_in[1]), 
        .grant(grant_1), .grant_v_o(grant_v[1]) );
  arbiter3_9 arbiter_w ( .clk(clk), .rst(rst), .request({\request[2][2] , 
        \request[2][1] , \request[2][0] }), .buffer_full_i(buffer_full_in[2]), 
        .grant(grant_2), .grant_v_o(grant_v[2]) );
  arbiter3_8 arbiter_l ( .clk(clk), .rst(rst), .request({\request[3][2] , 
        \request[3][1] , \request[3][0] }), .buffer_full_i(buffer_full_in[3]), 
        .grant(grant_3), .grant_v_o(grant_v[3]) );
  dccl_39 dccl_n ( .packet_addr_y_i({\packet_addr[0][3] , \packet_addr[0][2] , 
        \packet_addr[0][1] , \packet_addr[0][0] }), .packet_addr_x_i({
        \packet_addr[0][7] , \packet_addr[0][6] , \packet_addr[0][5] , 
        \packet_addr[0][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[0]), 
        .east_req(\request[1][0] ), .west_req(\request[2][0] ), .local_req(
        \request[3][0] ) );
  dccl_38 dccl_e ( .packet_addr_y_i({\packet_addr[1][3] , \packet_addr[1][2] , 
        \packet_addr[1][1] , \packet_addr[1][0] }), .packet_addr_x_i({
        \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] , 
        \packet_addr[1][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[1]), 
        .west_req(\request[2][1] ), .local_req(\request[3][1] ) );
  dccl_37 dccl_w ( .packet_addr_y_i({\packet_addr[2][3] , \packet_addr[2][2] , 
        \packet_addr[2][1] , \packet_addr[2][0] }), .packet_addr_x_i({
        \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] , 
        \packet_addr[2][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[2]), 
        .east_req(\request[1][1] ), .local_req(\request[3][2] ) );
  dccl_36 dccl_l ( .packet_addr_y_i({\packet_addr[3][3] , \packet_addr[3][2] , 
        \packet_addr[3][1] , \packet_addr[3][0] }), .packet_addr_x_i({
        \packet_addr[3][7] , \packet_addr[3][6] , \packet_addr[3][5] , 
        \packet_addr[3][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[3]), 
        .north_req(\request[0][0] ), .east_req(\request[1][2] ), .west_req(
        \request[2][2] ) );
endmodule


module mux3_1_10 ( data0, data1, data2, select0, select1, select2, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  output [15:0] data_o;
  input select0, select1, select2;
  wire   n1, n2, n6, n7, n8;

  AO222X1 U4 ( .IN1(data1[9]), .IN2(n8), .IN3(data0[9]), .IN4(n7), .IN5(
        data2[9]), .IN6(n6), .Q(data_o[9]) );
  AO222X1 U5 ( .IN1(data1[8]), .IN2(n8), .IN3(data0[8]), .IN4(n7), .IN5(
        data2[8]), .IN6(n6), .Q(data_o[8]) );
  AO222X1 U6 ( .IN1(data1[7]), .IN2(n8), .IN3(data0[7]), .IN4(n7), .IN5(
        data2[7]), .IN6(n6), .Q(data_o[7]) );
  AO222X1 U7 ( .IN1(data1[6]), .IN2(n8), .IN3(data0[6]), .IN4(n7), .IN5(
        data2[6]), .IN6(n6), .Q(data_o[6]) );
  AO222X1 U8 ( .IN1(data1[5]), .IN2(n8), .IN3(data0[5]), .IN4(n7), .IN5(
        data2[5]), .IN6(n6), .Q(data_o[5]) );
  AO222X1 U9 ( .IN1(data1[4]), .IN2(n8), .IN3(data0[4]), .IN4(n7), .IN5(
        data2[4]), .IN6(n6), .Q(data_o[4]) );
  AO222X1 U10 ( .IN1(data1[3]), .IN2(n8), .IN3(data0[3]), .IN4(n7), .IN5(
        data2[3]), .IN6(n6), .Q(data_o[3]) );
  AO222X1 U11 ( .IN1(data1[2]), .IN2(n8), .IN3(data0[2]), .IN4(n7), .IN5(
        data2[2]), .IN6(n6), .Q(data_o[2]) );
  AO222X1 U12 ( .IN1(data1[1]), .IN2(n8), .IN3(data0[1]), .IN4(n7), .IN5(
        data2[1]), .IN6(n6), .Q(data_o[1]) );
  AO222X1 U13 ( .IN1(data1[15]), .IN2(n8), .IN3(data0[15]), .IN4(n7), .IN5(
        data2[15]), .IN6(n6), .Q(data_o[15]) );
  AO222X1 U14 ( .IN1(data1[14]), .IN2(n8), .IN3(data0[14]), .IN4(n7), .IN5(
        data2[14]), .IN6(n6), .Q(data_o[14]) );
  AO222X1 U15 ( .IN1(data1[13]), .IN2(n8), .IN3(data0[13]), .IN4(n7), .IN5(
        data2[13]), .IN6(n6), .Q(data_o[13]) );
  AO222X1 U16 ( .IN1(data1[12]), .IN2(n8), .IN3(data0[12]), .IN4(n7), .IN5(
        data2[12]), .IN6(n6), .Q(data_o[12]) );
  AO222X1 U17 ( .IN1(data1[11]), .IN2(n8), .IN3(data0[11]), .IN4(n7), .IN5(
        data2[11]), .IN6(n6), .Q(data_o[11]) );
  AO222X1 U18 ( .IN1(data1[10]), .IN2(n8), .IN3(data0[10]), .IN4(n7), .IN5(
        data2[10]), .IN6(n6), .Q(data_o[10]) );
  AO222X1 U19 ( .IN1(data1[0]), .IN2(n8), .IN3(data0[0]), .IN4(n7), .IN5(
        data2[0]), .IN6(n6), .Q(data_o[0]) );
  INVX0 U2 ( .INP(select0), .ZN(n2) );
  INVX0 U3 ( .INP(select1), .ZN(n1) );
  AND3X1 U20 ( .IN1(n2), .IN2(n1), .IN3(select2), .Q(n6) );
  NOR3X0 U21 ( .IN1(select1), .IN2(select2), .IN3(n2), .QN(n7) );
  NOR3X0 U22 ( .IN1(select0), .IN2(select2), .IN3(n1), .QN(n8) );
endmodule


module mux3_1_9 ( data0, data1, data2, select0, select1, select2, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  output [15:0] data_o;
  input select0, select1, select2;
  wire   n1, n2, n6, n7, n8;

  AO222X1 U4 ( .IN1(data1[9]), .IN2(n8), .IN3(data0[9]), .IN4(n7), .IN5(
        data2[9]), .IN6(n6), .Q(data_o[9]) );
  AO222X1 U5 ( .IN1(data1[8]), .IN2(n8), .IN3(data0[8]), .IN4(n7), .IN5(
        data2[8]), .IN6(n6), .Q(data_o[8]) );
  AO222X1 U6 ( .IN1(data1[7]), .IN2(n8), .IN3(data0[7]), .IN4(n7), .IN5(
        data2[7]), .IN6(n6), .Q(data_o[7]) );
  AO222X1 U7 ( .IN1(data1[6]), .IN2(n8), .IN3(data0[6]), .IN4(n7), .IN5(
        data2[6]), .IN6(n6), .Q(data_o[6]) );
  AO222X1 U8 ( .IN1(data1[5]), .IN2(n8), .IN3(data0[5]), .IN4(n7), .IN5(
        data2[5]), .IN6(n6), .Q(data_o[5]) );
  AO222X1 U9 ( .IN1(data1[4]), .IN2(n8), .IN3(data0[4]), .IN4(n7), .IN5(
        data2[4]), .IN6(n6), .Q(data_o[4]) );
  AO222X1 U10 ( .IN1(data1[3]), .IN2(n8), .IN3(data0[3]), .IN4(n7), .IN5(
        data2[3]), .IN6(n6), .Q(data_o[3]) );
  AO222X1 U11 ( .IN1(data1[2]), .IN2(n8), .IN3(data0[2]), .IN4(n7), .IN5(
        data2[2]), .IN6(n6), .Q(data_o[2]) );
  AO222X1 U12 ( .IN1(data1[1]), .IN2(n8), .IN3(data0[1]), .IN4(n7), .IN5(
        data2[1]), .IN6(n6), .Q(data_o[1]) );
  AO222X1 U13 ( .IN1(data1[15]), .IN2(n8), .IN3(data0[15]), .IN4(n7), .IN5(
        data2[15]), .IN6(n6), .Q(data_o[15]) );
  AO222X1 U14 ( .IN1(data1[14]), .IN2(n8), .IN3(data0[14]), .IN4(n7), .IN5(
        data2[14]), .IN6(n6), .Q(data_o[14]) );
  AO222X1 U15 ( .IN1(data1[13]), .IN2(n8), .IN3(data0[13]), .IN4(n7), .IN5(
        data2[13]), .IN6(n6), .Q(data_o[13]) );
  AO222X1 U16 ( .IN1(data1[12]), .IN2(n8), .IN3(data0[12]), .IN4(n7), .IN5(
        data2[12]), .IN6(n6), .Q(data_o[12]) );
  AO222X1 U17 ( .IN1(data1[11]), .IN2(n8), .IN3(data0[11]), .IN4(n7), .IN5(
        data2[11]), .IN6(n6), .Q(data_o[11]) );
  AO222X1 U18 ( .IN1(data1[10]), .IN2(n8), .IN3(data0[10]), .IN4(n7), .IN5(
        data2[10]), .IN6(n6), .Q(data_o[10]) );
  AO222X1 U19 ( .IN1(data1[0]), .IN2(n8), .IN3(data0[0]), .IN4(n7), .IN5(
        data2[0]), .IN6(n6), .Q(data_o[0]) );
  INVX0 U2 ( .INP(select0), .ZN(n2) );
  INVX0 U3 ( .INP(select1), .ZN(n1) );
  AND3X1 U20 ( .IN1(n2), .IN2(n1), .IN3(select2), .Q(n6) );
  NOR3X0 U21 ( .IN1(select1), .IN2(select2), .IN3(n2), .QN(n7) );
  NOR3X0 U22 ( .IN1(select0), .IN2(select2), .IN3(n1), .QN(n8) );
endmodule


module mux3_1_8 ( data0, data1, data2, select0, select1, select2, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  output [15:0] data_o;
  input select0, select1, select2;
  wire   n1, n2, n6, n7, n8;

  AO222X1 U4 ( .IN1(data1[9]), .IN2(n8), .IN3(data0[9]), .IN4(n7), .IN5(
        data2[9]), .IN6(n6), .Q(data_o[9]) );
  AO222X1 U5 ( .IN1(data1[8]), .IN2(n8), .IN3(data0[8]), .IN4(n7), .IN5(
        data2[8]), .IN6(n6), .Q(data_o[8]) );
  AO222X1 U6 ( .IN1(data1[7]), .IN2(n8), .IN3(data0[7]), .IN4(n7), .IN5(
        data2[7]), .IN6(n6), .Q(data_o[7]) );
  AO222X1 U7 ( .IN1(data1[6]), .IN2(n8), .IN3(data0[6]), .IN4(n7), .IN5(
        data2[6]), .IN6(n6), .Q(data_o[6]) );
  AO222X1 U8 ( .IN1(data1[5]), .IN2(n8), .IN3(data0[5]), .IN4(n7), .IN5(
        data2[5]), .IN6(n6), .Q(data_o[5]) );
  AO222X1 U9 ( .IN1(data1[4]), .IN2(n8), .IN3(data0[4]), .IN4(n7), .IN5(
        data2[4]), .IN6(n6), .Q(data_o[4]) );
  AO222X1 U10 ( .IN1(data1[3]), .IN2(n8), .IN3(data0[3]), .IN4(n7), .IN5(
        data2[3]), .IN6(n6), .Q(data_o[3]) );
  AO222X1 U11 ( .IN1(data1[2]), .IN2(n8), .IN3(data0[2]), .IN4(n7), .IN5(
        data2[2]), .IN6(n6), .Q(data_o[2]) );
  AO222X1 U12 ( .IN1(data1[1]), .IN2(n8), .IN3(data0[1]), .IN4(n7), .IN5(
        data2[1]), .IN6(n6), .Q(data_o[1]) );
  AO222X1 U13 ( .IN1(data1[15]), .IN2(n8), .IN3(data0[15]), .IN4(n7), .IN5(
        data2[15]), .IN6(n6), .Q(data_o[15]) );
  AO222X1 U14 ( .IN1(data1[14]), .IN2(n8), .IN3(data0[14]), .IN4(n7), .IN5(
        data2[14]), .IN6(n6), .Q(data_o[14]) );
  AO222X1 U15 ( .IN1(data1[13]), .IN2(n8), .IN3(data0[13]), .IN4(n7), .IN5(
        data2[13]), .IN6(n6), .Q(data_o[13]) );
  AO222X1 U16 ( .IN1(data1[12]), .IN2(n8), .IN3(data0[12]), .IN4(n7), .IN5(
        data2[12]), .IN6(n6), .Q(data_o[12]) );
  AO222X1 U17 ( .IN1(data1[11]), .IN2(n8), .IN3(data0[11]), .IN4(n7), .IN5(
        data2[11]), .IN6(n6), .Q(data_o[11]) );
  AO222X1 U18 ( .IN1(data1[10]), .IN2(n8), .IN3(data0[10]), .IN4(n7), .IN5(
        data2[10]), .IN6(n6), .Q(data_o[10]) );
  AO222X1 U19 ( .IN1(data1[0]), .IN2(n8), .IN3(data0[0]), .IN4(n7), .IN5(
        data2[0]), .IN6(n6), .Q(data_o[0]) );
  INVX0 U2 ( .INP(select0), .ZN(n2) );
  INVX0 U3 ( .INP(select1), .ZN(n1) );
  AND3X1 U20 ( .IN1(n2), .IN2(n1), .IN3(select2), .Q(n6) );
  NOR3X0 U21 ( .IN1(select1), .IN2(select2), .IN3(n2), .QN(n7) );
  NOR3X0 U22 ( .IN1(select0), .IN2(select2), .IN3(n1), .QN(n8) );
endmodule



    module node4_NODE_X2_NODE_Y3I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__I_node_2_node_interface__ ( 
        \clk.clk , \reset.reset , \local_node.clk , 
        \local_node.buffer_full_in , \local_node.buffer_full_out , 
        \local_node.receiving_data , \local_node.sending_data , 
        \local_node.data_in , \local_node.data_out , \node_0.clk , 
        \node_0.buffer_full_in , \node_0.buffer_full_out , 
        \node_0.receiving_data , \node_0.sending_data , \node_0.data_in , 
        \node_0.data_out , \node_1.clk , \node_1.buffer_full_in , 
        \node_1.buffer_full_out , \node_1.receiving_data , 
        \node_1.sending_data , \node_1.data_in , \node_1.data_out , 
        \node_2.clk , \node_2.buffer_full_in , \node_2.buffer_full_out , 
        \node_2.receiving_data , \node_2.sending_data , \node_2.data_in , 
        \node_2.data_out  );
  input [15:0] \local_node.data_in ;
  output [15:0] \local_node.data_out ;
  input [15:0] \node_0.data_in ;
  output [15:0] \node_0.data_out ;
  input [15:0] \node_1.data_in ;
  output [15:0] \node_1.data_out ;
  input [15:0] \node_2.data_in ;
  output [15:0] \node_2.data_out ;
  input \clk.clk , \reset.reset , \local_node.buffer_full_in ,
         \local_node.receiving_data , \node_0.buffer_full_in ,
         \node_0.receiving_data , \node_1.buffer_full_in ,
         \node_1.receiving_data , \node_2.buffer_full_in ,
         \node_2.receiving_data ;
  output \local_node.buffer_full_out , \local_node.sending_data ,
         \node_0.buffer_full_out , \node_0.sending_data ,
         \node_1.buffer_full_out , \node_1.sending_data ,
         \node_2.buffer_full_out , \node_2.sending_data ;
  inout \local_node.clk ,  \node_0.clk ,  \node_1.clk ,  \node_2.clk ;
  wire   \buffer_out[3][15] , \buffer_out[3][14] , \buffer_out[3][13] ,
         \buffer_out[3][12] , \buffer_out[3][11] , \buffer_out[3][10] ,
         \buffer_out[3][9] , \buffer_out[3][8] , \buffer_out[3][7] ,
         \buffer_out[3][6] , \buffer_out[3][5] , \buffer_out[3][4] ,
         \buffer_out[3][3] , \buffer_out[3][2] , \buffer_out[3][1] ,
         \buffer_out[3][0] , \buffer_out[2][15] , \buffer_out[2][14] ,
         \buffer_out[2][13] , \buffer_out[2][12] , \buffer_out[2][11] ,
         \buffer_out[2][10] , \buffer_out[2][9] , \buffer_out[2][8] ,
         \buffer_out[2][7] , \buffer_out[2][6] , \buffer_out[2][5] ,
         \buffer_out[2][4] , \buffer_out[2][3] , \buffer_out[2][2] ,
         \buffer_out[2][1] , \buffer_out[2][0] , \buffer_out[1][15] ,
         \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] ,
         \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] ,
         \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] ,
         \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] ,
         \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] ,
         \buffer_out[0][15] , \buffer_out[0][14] , \buffer_out[0][13] ,
         \buffer_out[0][12] , \buffer_out[0][11] , \buffer_out[0][10] ,
         \buffer_out[0][9] , \buffer_out[0][8] , \buffer_out[0][7] ,
         \buffer_out[0][6] , \buffer_out[0][5] , \buffer_out[0][4] ,
         \buffer_out[0][3] , \buffer_out[0][2] , \buffer_out[0][1] ,
         \buffer_out[0][0] , \next_buffer_out[3][15] ,
         \next_buffer_out[3][14] , \next_buffer_out[3][13] ,
         \next_buffer_out[3][12] , \next_buffer_out[3][11] ,
         \next_buffer_out[3][10] , \next_buffer_out[3][9] ,
         \next_buffer_out[3][8] , \next_buffer_out[3][7] ,
         \next_buffer_out[3][6] , \next_buffer_out[3][5] ,
         \next_buffer_out[3][4] , \next_buffer_out[3][3] ,
         \next_buffer_out[3][2] , \next_buffer_out[3][1] ,
         \next_buffer_out[3][0] , \next_buffer_out[2][15] ,
         \next_buffer_out[2][14] , \next_buffer_out[2][13] ,
         \next_buffer_out[2][12] , \next_buffer_out[2][11] ,
         \next_buffer_out[2][10] , \next_buffer_out[2][9] ,
         \next_buffer_out[2][8] , \next_buffer_out[2][7] ,
         \next_buffer_out[2][6] , \next_buffer_out[2][5] ,
         \next_buffer_out[2][4] , \next_buffer_out[2][3] ,
         \next_buffer_out[2][2] , \next_buffer_out[2][1] ,
         \next_buffer_out[2][0] , \next_buffer_out[1][15] ,
         \next_buffer_out[1][14] , \next_buffer_out[1][13] ,
         \next_buffer_out[1][12] , \next_buffer_out[1][11] ,
         \next_buffer_out[1][10] , \next_buffer_out[1][9] ,
         \next_buffer_out[1][8] , \next_buffer_out[1][7] ,
         \next_buffer_out[1][6] , \next_buffer_out[1][5] ,
         \next_buffer_out[1][4] , \next_buffer_out[1][3] ,
         \next_buffer_out[1][2] , \next_buffer_out[1][1] ,
         \next_buffer_out[1][0] , \next_buffer_out[0][15] ,
         \next_buffer_out[0][14] , \next_buffer_out[0][13] ,
         \next_buffer_out[0][12] , \next_buffer_out[0][11] ,
         \next_buffer_out[0][10] , \next_buffer_out[0][9] ,
         \next_buffer_out[0][8] , \next_buffer_out[0][7] ,
         \next_buffer_out[0][6] , \next_buffer_out[0][5] ,
         \next_buffer_out[0][4] , \next_buffer_out[0][3] ,
         \next_buffer_out[0][2] , \next_buffer_out[0][1] ,
         \next_buffer_out[0][0] ;
  wire   [3:0] buffer_full_in;
  wire   [3:0] receiving_data;
  wire   [3:0] pop_v;
  wire   [3:0] data_valid;
  wire   [3:0] next_data_valid;
  wire   [2:0] grant_1;
  wire   [2:0] grant_2;
  wire   [2:0] grant_3;
  tri   \local_node.buffer_full_in ;
  tri   \local_node.buffer_full_out ;
  tri   \local_node.receiving_data ;
  tri   \local_node.sending_data ;
  tri   [15:0] \local_node.data_in ;
  tri   [15:0] \local_node.data_out ;

  converter_out_I_n_node_interface_dut_ c3 ( .\n.buffer_full_in (
        \local_node.buffer_full_in ), .\n.receiving_data (
        \local_node.receiving_data ), .\n.data_in (\local_node.data_in ), 
        .\n.buffer_full_out (\local_node.buffer_full_out ), .\n.sending_data (
        \local_node.sending_data ), .\n.data_out (\local_node.data_out ), 
        .buffer_full_in(1'b0), .receiving_data(1'b0), .data_in({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  fifo_kev_39 \genblk1[0].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[0]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[0]), .data_out({\buffer_out[0][15] , 
        \buffer_out[0][14] , \buffer_out[0][13] , \buffer_out[0][12] , 
        \buffer_out[0][11] , \buffer_out[0][10] , \buffer_out[0][9] , 
        \buffer_out[0][8] , \buffer_out[0][7] , \buffer_out[0][6] , 
        \buffer_out[0][5] , \buffer_out[0][4] , \buffer_out[0][3] , 
        \buffer_out[0][2] , \buffer_out[0][1] , \buffer_out[0][0] }), 
        .next_data_out({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] , 
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .next_data_valid(
        next_data_valid[0]) );
  address_counter_39 \genblk1[0].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] }), 
        .buffer_data_valid(next_data_valid[0]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .buffer_pop(
        pop_v[0]), .receiving_data(1'b0) );
  fifo_kev_38 \genblk1[1].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[1]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[1]), .data_out({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), 
        .next_data_out({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] , 
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .next_data_valid(
        next_data_valid[1]) );
  address_counter_38 \genblk1[1].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] }), 
        .buffer_data_valid(next_data_valid[1]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .buffer_pop(
        pop_v[1]), .receiving_data(1'b0) );
  fifo_kev_37 \genblk1[2].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[2]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[2]), .data_out({\buffer_out[2][15] , 
        \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] , 
        \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] , 
        \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] , 
        \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] , 
        \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] }), 
        .next_data_out({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] , 
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .next_data_valid(
        next_data_valid[2]) );
  address_counter_37 \genblk1[2].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] }), 
        .buffer_data_valid(next_data_valid[2]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .buffer_pop(
        pop_v[2]), .receiving_data(1'b0) );
  fifo_kev_36 \genblk1[3].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[3]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[3]), .data_out({\buffer_out[3][15] , 
        \buffer_out[3][14] , \buffer_out[3][13] , \buffer_out[3][12] , 
        \buffer_out[3][11] , \buffer_out[3][10] , \buffer_out[3][9] , 
        \buffer_out[3][8] , \buffer_out[3][7] , \buffer_out[3][6] , 
        \buffer_out[3][5] , \buffer_out[3][4] , \buffer_out[3][3] , 
        \buffer_out[3][2] , \buffer_out[3][1] , \buffer_out[3][0] }), 
        .next_data_out({\next_buffer_out[3][15] , \next_buffer_out[3][14] , 
        \next_buffer_out[3][13] , \next_buffer_out[3][12] , 
        \next_buffer_out[3][11] , \next_buffer_out[3][10] , 
        \next_buffer_out[3][9] , \next_buffer_out[3][8] , 
        \next_buffer_out[3][7] , \next_buffer_out[3][6] , 
        \next_buffer_out[3][5] , \next_buffer_out[3][4] , 
        \next_buffer_out[3][3] , \next_buffer_out[3][2] , 
        \next_buffer_out[3][1] , \next_buffer_out[3][0] }), .next_data_valid(
        next_data_valid[3]) );
  address_counter_36 \genblk1[3].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[3][15] , \next_buffer_out[3][14] , 
        \next_buffer_out[3][13] , \next_buffer_out[3][12] , 
        \next_buffer_out[3][11] , \next_buffer_out[3][10] , 
        \next_buffer_out[3][9] , \next_buffer_out[3][8] }), 
        .buffer_data_valid(next_data_valid[3]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[3][7] , \next_buffer_out[3][6] , 
        \next_buffer_out[3][5] , \next_buffer_out[3][4] , 
        \next_buffer_out[3][3] , \next_buffer_out[3][2] , 
        \next_buffer_out[3][1] , \next_buffer_out[3][0] }), .buffer_pop(
        pop_v[3]), .receiving_data(1'b0) );
  converter_in_I_n_node_interface_dut__15 \genblk2.c0  ( .\n.buffer_full_in (
        \node_0.buffer_full_in ), .\n.receiving_data (\node_0.receiving_data ), 
        .\n.data_in (\node_0.data_in ), .\n.buffer_full_out (
        \node_0.buffer_full_out ), .\n.sending_data (\node_0.sending_data ), 
        .\n.data_out (\node_0.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_in_I_n_node_interface_dut__14 \genblk2.c1  ( .\n.buffer_full_in (
        \node_1.buffer_full_in ), .\n.receiving_data (\node_1.receiving_data ), 
        .\n.data_in (\node_1.data_in ), .\n.buffer_full_out (
        \node_1.buffer_full_out ), .\n.sending_data (\node_1.sending_data ), 
        .\n.data_out (\node_1.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_out_I_n_node_interface_dut_ \genblk2.c2  ( .\n.buffer_full_in (
        \node_2.buffer_full_in ), .\n.receiving_data (\node_2.receiving_data ), 
        .\n.data_in (\node_2.data_in ), .\n.buffer_full_out (
        \node_2.buffer_full_out ), .\n.sending_data (\node_2.sending_data ), 
        .\n.data_out (\node_2.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  controller4_edge_s_0 \genblk2.s  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .packet_addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .local_addr({1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1}), 
        .packet_valid(data_valid), .buffer_full_in({1'b0, 1'b0, 1'b0, 1'b0}), 
        .grant_1(grant_1), .grant_2(grant_2), .grant_3(grant_3), .pop_v(pop_v)
         );
  mux3_1_10 \genblk2.mux_e  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[2][15] , 
        \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] , 
        \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] , 
        \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] , 
        \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] , 
        \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] }), .data2({
        \buffer_out[3][15] , \buffer_out[3][14] , \buffer_out[3][13] , 
        \buffer_out[3][12] , \buffer_out[3][11] , \buffer_out[3][10] , 
        \buffer_out[3][9] , \buffer_out[3][8] , \buffer_out[3][7] , 
        \buffer_out[3][6] , \buffer_out[3][5] , \buffer_out[3][4] , 
        \buffer_out[3][3] , \buffer_out[3][2] , \buffer_out[3][1] , 
        \buffer_out[3][0] }), .select0(grant_1[0]), .select1(grant_1[1]), 
        .select2(grant_1[2]) );
  mux3_1_9 \genblk2.mux_w  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[3][15] , \buffer_out[3][14] , \buffer_out[3][13] , 
        \buffer_out[3][12] , \buffer_out[3][11] , \buffer_out[3][10] , 
        \buffer_out[3][9] , \buffer_out[3][8] , \buffer_out[3][7] , 
        \buffer_out[3][6] , \buffer_out[3][5] , \buffer_out[3][4] , 
        \buffer_out[3][3] , \buffer_out[3][2] , \buffer_out[3][1] , 
        \buffer_out[3][0] }), .select0(grant_2[0]), .select1(grant_2[1]), 
        .select2(grant_2[2]) );
  mux3_1_8 \genblk2.mux_l  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[2][15] , \buffer_out[2][14] , \buffer_out[2][13] , 
        \buffer_out[2][12] , \buffer_out[2][11] , \buffer_out[2][10] , 
        \buffer_out[2][9] , \buffer_out[2][8] , \buffer_out[2][7] , 
        \buffer_out[2][6] , \buffer_out[2][5] , \buffer_out[2][4] , 
        \buffer_out[2][3] , \buffer_out[2][2] , \buffer_out[2][1] , 
        \buffer_out[2][0] }), .select0(grant_3[0]), .select1(grant_3[1]), 
        .select2(grant_3[2]) );
endmodule


module fifo_kev_35 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_71 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_35 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_71 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_70 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_35 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_70 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_35_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_35 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_35 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_35 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_35_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_34 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_69 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_34 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_69 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_68 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_34 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_68 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_34_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_34 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_34 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_34 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_34_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_33 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_67 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_33 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_67 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_66 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_33 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_66 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_33_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_33 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_33 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_33 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_33_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_32 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_65 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_32 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_65 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_64 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_32 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_64 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_32_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_32 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_32 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_32 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_32_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module converter_in_I_n_node_interface_dut__13 ( \n.buffer_full_in , 
        \n.receiving_data , \n.data_in , \n.buffer_full_out , \n.sending_data , 
        \n.data_out , buffer_full_out, sending_data, data_out, buffer_full_in, 
        receiving_data, data_in );
  input [15:0] \n.data_in ;
  output [15:0] \n.data_out ;
  output [15:0] data_out;
  input [15:0] data_in;
  input \n.buffer_full_in , \n.receiving_data , buffer_full_in, receiving_data;
  output \n.buffer_full_out , \n.sending_data , buffer_full_out, sending_data;
  wire   \n.buffer_full_in , \n.receiving_data , buffer_full_in,
         receiving_data;
  assign buffer_full_out = \n.buffer_full_in ;
  assign sending_data = \n.receiving_data ;
  assign data_out[15] = \n.data_in  [15];
  assign data_out[14] = \n.data_in  [14];
  assign data_out[13] = \n.data_in  [13];
  assign data_out[12] = \n.data_in  [12];
  assign data_out[11] = \n.data_in  [11];
  assign data_out[10] = \n.data_in  [10];
  assign data_out[9] = \n.data_in  [9];
  assign data_out[8] = \n.data_in  [8];
  assign data_out[7] = \n.data_in  [7];
  assign data_out[6] = \n.data_in  [6];
  assign data_out[5] = \n.data_in  [5];
  assign data_out[4] = \n.data_in  [4];
  assign data_out[3] = \n.data_in  [3];
  assign data_out[2] = \n.data_in  [2];
  assign data_out[1] = \n.data_in  [1];
  assign data_out[0] = \n.data_in  [0];
  assign \n.buffer_full_out  = buffer_full_in;
  assign \n.sending_data  = receiving_data;
  assign \n.data_out  [15] = data_in[15];
  assign \n.data_out  [14] = data_in[14];
  assign \n.data_out  [13] = data_in[13];
  assign \n.data_out  [12] = data_in[12];
  assign \n.data_out  [11] = data_in[11];
  assign \n.data_out  [10] = data_in[10];
  assign \n.data_out  [9] = data_in[9];
  assign \n.data_out  [8] = data_in[8];
  assign \n.data_out  [7] = data_in[7];
  assign \n.data_out  [6] = data_in[6];
  assign \n.data_out  [5] = data_in[5];
  assign \n.data_out  [4] = data_in[4];
  assign \n.data_out  [3] = data_in[3];
  assign \n.data_out  [2] = data_in[2];
  assign \n.data_out  [1] = data_in[1];
  assign \n.data_out  [0] = data_in[0];

endmodule


module converter_in_I_n_node_interface_dut__12 ( \n.buffer_full_in , 
        \n.receiving_data , \n.data_in , \n.buffer_full_out , \n.sending_data , 
        \n.data_out , buffer_full_out, sending_data, data_out, buffer_full_in, 
        receiving_data, data_in );
  input [15:0] \n.data_in ;
  output [15:0] \n.data_out ;
  output [15:0] data_out;
  input [15:0] data_in;
  input \n.buffer_full_in , \n.receiving_data , buffer_full_in, receiving_data;
  output \n.buffer_full_out , \n.sending_data , buffer_full_out, sending_data;
  wire   \n.buffer_full_in , \n.receiving_data , buffer_full_in,
         receiving_data;
  assign buffer_full_out = \n.buffer_full_in ;
  assign sending_data = \n.receiving_data ;
  assign data_out[15] = \n.data_in  [15];
  assign data_out[14] = \n.data_in  [14];
  assign data_out[13] = \n.data_in  [13];
  assign data_out[12] = \n.data_in  [12];
  assign data_out[11] = \n.data_in  [11];
  assign data_out[10] = \n.data_in  [10];
  assign data_out[9] = \n.data_in  [9];
  assign data_out[8] = \n.data_in  [8];
  assign data_out[7] = \n.data_in  [7];
  assign data_out[6] = \n.data_in  [6];
  assign data_out[5] = \n.data_in  [5];
  assign data_out[4] = \n.data_in  [4];
  assign data_out[3] = \n.data_in  [3];
  assign data_out[2] = \n.data_in  [2];
  assign data_out[1] = \n.data_in  [1];
  assign data_out[0] = \n.data_in  [0];
  assign \n.buffer_full_out  = buffer_full_in;
  assign \n.sending_data  = receiving_data;
  assign \n.data_out  [15] = data_in[15];
  assign \n.data_out  [14] = data_in[14];
  assign \n.data_out  [13] = data_in[13];
  assign \n.data_out  [12] = data_in[12];
  assign \n.data_out  [11] = data_in[11];
  assign \n.data_out  [10] = data_in[10];
  assign \n.data_out  [9] = data_in[9];
  assign \n.data_out  [8] = data_in[8];
  assign \n.data_out  [7] = data_in[7];
  assign \n.data_out  [6] = data_in[6];
  assign \n.data_out  [5] = data_in[5];
  assign \n.data_out  [4] = data_in[4];
  assign \n.data_out  [3] = data_in[3];
  assign \n.data_out  [2] = data_in[2];
  assign \n.data_out  [1] = data_in[1];
  assign \n.data_out  [0] = data_in[0];

endmodule


module flipflop_BITS2_15 ( clk, data_i, data_o );
  input [1:0] data_i;
  output [1:0] data_o;
  input clk;


  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS2_15 ( clk, enable_i, reset, data_i, data_o );
  input [1:0] data_i;
  input [1:0] data_o;
  input clk, enable_i, reset;
  wire   n10, n11, n1, n5, n7, n8, n9;
  wire   [1:0] write_data;

  AOI22X1 U5 ( .IN1(enable_i), .IN2(data_i[1]), .IN3(n10), .IN4(n1), .QN(n9)
         );
  AOI22X1 U6 ( .IN1(data_i[0]), .IN2(enable_i), .IN3(n11), .IN4(n1), .QN(n8)
         );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n9), .QN(write_data[1]) );
  NOR2X0 U4 ( .IN1(reset), .IN2(n8), .QN(write_data[0]) );
  AND2X1 U7 ( .IN1(data_o[1]), .IN2(n7), .Q(n10) );
  AND2X1 U8 ( .IN1(data_o[0]), .IN2(n5), .Q(n11) );
  flipflop_BITS2_15 FF ( .clk(clk), .data_i(write_data), .data_o({n7, n5}) );
endmodule


module flipflop_BITS1_55 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_55 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_55 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter2_15 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [1:0] request;
  output [1:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   tail_en, n1, n2;
  wire   [1:0] req_i;
  wire   [1:0] req_o;

  AND3X1 U10 ( .IN1(request[1]), .IN2(n1), .IN3(n2), .Q(grant[1]) );
  AND3X1 U11 ( .IN1(request[0]), .IN2(n2), .IN3(request[1]), .Q(tail_en) );
  INVX0 U6 ( .INP(request[0]), .ZN(n1) );
  NOR2X0 U7 ( .IN1(buffer_full_i), .IN2(n1), .QN(grant[0]) );
  INVX0 U8 ( .INP(buffer_full_i), .ZN(n2) );
  OA21X1 U9 ( .IN1(request[1]), .IN2(request[0]), .IN3(n2), .Q(grant_v_o) );
  register_BITS2_15 req_record ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i({1'b1, 1'b0}), .data_o({1'b0, 1'b0}) );
  register_BITS1_55 tail ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i(1'b1), .data_o(1'b0) );
endmodule


module flipflop_BITS2_14 ( clk, data_i, data_o );
  input [1:0] data_i;
  output [1:0] data_o;
  input clk;


  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS2_14 ( clk, enable_i, reset, data_i, data_o );
  input [1:0] data_i;
  input [1:0] data_o;
  input clk, enable_i, reset;
  wire   n10, n11, n1, n5, n7, n8, n9;
  wire   [1:0] write_data;

  AOI22X1 U5 ( .IN1(enable_i), .IN2(data_i[1]), .IN3(n10), .IN4(n1), .QN(n9)
         );
  AOI22X1 U6 ( .IN1(data_i[0]), .IN2(enable_i), .IN3(n11), .IN4(n1), .QN(n8)
         );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n9), .QN(write_data[1]) );
  NOR2X0 U4 ( .IN1(reset), .IN2(n8), .QN(write_data[0]) );
  AND2X1 U7 ( .IN1(data_o[1]), .IN2(n7), .Q(n10) );
  AND2X1 U8 ( .IN1(data_o[0]), .IN2(n5), .Q(n11) );
  flipflop_BITS2_14 FF ( .clk(clk), .data_i(write_data), .data_o({n7, n5}) );
endmodule


module flipflop_BITS1_54 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_54 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_54 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter2_14 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [1:0] request;
  output [1:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   tail_en, n1, n2;
  wire   [1:0] req_i;
  wire   [1:0] req_o;

  AND3X1 U10 ( .IN1(request[1]), .IN2(n1), .IN3(n2), .Q(grant[1]) );
  AND3X1 U11 ( .IN1(request[0]), .IN2(n2), .IN3(request[1]), .Q(tail_en) );
  INVX0 U6 ( .INP(request[0]), .ZN(n1) );
  NOR2X0 U7 ( .IN1(buffer_full_i), .IN2(n1), .QN(grant[0]) );
  INVX0 U8 ( .INP(buffer_full_i), .ZN(n2) );
  OA21X1 U9 ( .IN1(request[1]), .IN2(request[0]), .IN3(n2), .Q(grant_v_o) );
  register_BITS2_14 req_record ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i({1'b1, 1'b0}), .data_o({1'b0, 1'b0}) );
  register_BITS1_54 tail ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i(1'b1), .data_o(1'b0) );
endmodule


module flipflop_BITS3_15 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_15 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_15 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS3_14 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_14 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_14 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS1_53 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_53 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_53 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_52 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_52 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_52 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter3_7 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [2:0] request;
  output [2:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[1][2] , \req_i[1][1] , \req_i[1][0] , \req_i[0][2] ,
         \req_i[0][1] , tail_en, N99, N100, N101, N110, N111, N118, N119, N120,
         N121, n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [1:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N99 = request[0];
  assign N100 = request[1];
  assign N101 = request[2];

  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(N111), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(N110), .Q(\req_i[0][1] ) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N121), .D(tail_en), .Q(req_en[0]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N120), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N119), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N118), .Q(grant[0]) );
  AND2X1 U20 ( .IN1(n8), .IN2(N101), .Q(n7) );
  OR3X1 U21 ( .IN1(n3), .IN2(N111), .IN3(n6), .Q(N121) );
  NOR3X0 U22 ( .IN1(N99), .IN2(N100), .IN3(n6), .QN(N120) );
  NOR3X0 U23 ( .IN1(n2), .IN2(N99), .IN3(n6), .QN(N119) );
  NAND3X0 U24 ( .IN1(n2), .IN2(n3), .IN3(n1), .QN(n5) );
  AO22X1 U25 ( .IN1(N100), .IN2(N101), .IN3(N99), .IN4(N101), .Q(N111) );
  INVX0 U10 ( .INP(N101), .ZN(n3) );
  NAND2X1 U11 ( .IN1(n5), .IN2(n4), .QN(n6) );
  INVX0 U12 ( .INP(N99), .ZN(n1) );
  INVX0 U13 ( .INP(N100), .ZN(n2) );
  INVX0 U14 ( .INP(buffer_full_i), .ZN(n4) );
  NAND2X1 U15 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NOR2X0 U16 ( .IN1(n1), .IN2(n6), .QN(N118) );
  NOR2X0 U17 ( .IN1(n1), .IN2(n2), .QN(N110) );
  OA21X1 U18 ( .IN1(N110), .IN2(n7), .IN3(n4), .Q(tail_en) );
  OA21X1 U19 ( .IN1(N101), .IN2(n8), .IN3(n4), .Q(grant_v_o) );
  register_BITS3_15 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][2] , \req_i[0][1] , 1'b0}), .data_o({
        1'b0, 1'b0, 1'b0}) );
  register_BITS3_14 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][2] , \req_i[1][1] , \req_i[1][0] }), 
        .data_o({1'b0, 1'b0, 1'b0}) );
  register_BITS1_53 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b1), .data_o(1'b0) );
  register_BITS1_52 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module flipflop_BITS3_13 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_13 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_13 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS3_12 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_12 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_12 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS1_51 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_51 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_51 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_50 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_50 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_50 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter3_6 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [2:0] request;
  output [2:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[1][2] , \req_i[1][1] , \req_i[1][0] , \req_i[0][2] ,
         \req_i[0][1] , tail_en, N99, N100, N101, N110, N111, N118, N119, N120,
         N121, n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [1:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N99 = request[0];
  assign N100 = request[1];
  assign N101 = request[2];

  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(N111), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(N110), .Q(\req_i[0][1] ) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N121), .D(tail_en), .Q(req_en[0]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N120), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N119), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N118), .Q(grant[0]) );
  AND2X1 U20 ( .IN1(n8), .IN2(N101), .Q(n7) );
  OR3X1 U21 ( .IN1(n3), .IN2(N111), .IN3(n6), .Q(N121) );
  NOR3X0 U22 ( .IN1(N99), .IN2(N100), .IN3(n6), .QN(N120) );
  NOR3X0 U23 ( .IN1(n2), .IN2(N99), .IN3(n6), .QN(N119) );
  NAND3X0 U24 ( .IN1(n2), .IN2(n3), .IN3(n1), .QN(n5) );
  AO22X1 U25 ( .IN1(N100), .IN2(N101), .IN3(N99), .IN4(N101), .Q(N111) );
  INVX0 U10 ( .INP(N101), .ZN(n3) );
  NAND2X1 U11 ( .IN1(n5), .IN2(n4), .QN(n6) );
  INVX0 U12 ( .INP(N99), .ZN(n1) );
  INVX0 U13 ( .INP(N100), .ZN(n2) );
  INVX0 U14 ( .INP(buffer_full_i), .ZN(n4) );
  NAND2X1 U15 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NOR2X0 U16 ( .IN1(n1), .IN2(n6), .QN(N118) );
  NOR2X0 U17 ( .IN1(n1), .IN2(n2), .QN(N110) );
  OA21X1 U18 ( .IN1(N110), .IN2(n7), .IN3(n4), .Q(tail_en) );
  OA21X1 U19 ( .IN1(N101), .IN2(n8), .IN3(n4), .Q(grant_v_o) );
  register_BITS3_13 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][2] , \req_i[0][1] , 1'b0}), .data_o({
        1'b0, 1'b0, 1'b0}) );
  register_BITS3_12 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][2] , \req_i[1][1] , \req_i[1][0] }), 
        .data_o({1'b0, 1'b0, 1'b0}) );
  register_BITS1_51 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b1), .data_o(1'b0) );
  register_BITS1_50 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module dccl_35 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_34 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_33 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_32 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module controller4_edge_w_1 ( clk, rst, .packet_addr({\packet_addr[3][7] , 
        \packet_addr[3][6] , \packet_addr[3][5] , \packet_addr[3][4] , 
        \packet_addr[3][3] , \packet_addr[3][2] , \packet_addr[3][1] , 
        \packet_addr[3][0] , \packet_addr[2][7] , \packet_addr[2][6] , 
        \packet_addr[2][5] , \packet_addr[2][4] , \packet_addr[2][3] , 
        \packet_addr[2][2] , \packet_addr[2][1] , \packet_addr[2][0] , 
        \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] , 
        \packet_addr[1][4] , \packet_addr[1][3] , \packet_addr[1][2] , 
        \packet_addr[1][1] , \packet_addr[1][0] , \packet_addr[0][7] , 
        \packet_addr[0][6] , \packet_addr[0][5] , \packet_addr[0][4] , 
        \packet_addr[0][3] , \packet_addr[0][2] , \packet_addr[0][1] , 
        \packet_addr[0][0] }), local_addr, packet_valid, buffer_full_in, 
        grant_0, grant_1, grant_2, grant_3, grant_v, pop_v );
  input [7:0] local_addr;
  input [3:0] packet_valid;
  input [3:0] buffer_full_in;
  output [1:0] grant_0;
  output [1:0] grant_1;
  output [2:0] grant_2;
  output [2:0] grant_3;
  output [3:0] grant_v;
  output [3:0] pop_v;
  input clk, rst, \packet_addr[3][7] , \packet_addr[3][6] ,
         \packet_addr[3][5] , \packet_addr[3][4] , \packet_addr[3][3] ,
         \packet_addr[3][2] , \packet_addr[3][1] , \packet_addr[3][0] ,
         \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] ,
         \packet_addr[2][4] , \packet_addr[2][3] , \packet_addr[2][2] ,
         \packet_addr[2][1] , \packet_addr[2][0] , \packet_addr[1][7] ,
         \packet_addr[1][6] , \packet_addr[1][5] , \packet_addr[1][4] ,
         \packet_addr[1][3] , \packet_addr[1][2] , \packet_addr[1][1] ,
         \packet_addr[1][0] , \packet_addr[0][7] , \packet_addr[0][6] ,
         \packet_addr[0][5] , \packet_addr[0][4] , \packet_addr[0][3] ,
         \packet_addr[0][2] , \packet_addr[0][1] , \packet_addr[0][0] ;
  wire   \grant_3[2] , \request[3][2] , \request[3][1] , \request[3][0] ,
         \request[2][2] , \request[2][1] , \request[2][0] , \request[1][1] ,
         \request[1][0] , \request[0][1] , \request[0][0] ;
  assign pop_v[2] = \grant_3[2] ;
  assign grant_3[2] = \grant_3[2] ;

  OR3X1 U1 ( .IN1(grant_2[2]), .IN2(grant_1[1]), .IN3(grant_0[1]), .Q(pop_v[3]) );
  OR3X1 U2 ( .IN1(grant_3[1]), .IN2(grant_2[1]), .IN3(grant_0[0]), .Q(pop_v[1]) );
  OR3X1 U3 ( .IN1(grant_3[0]), .IN2(grant_2[0]), .IN3(grant_1[0]), .Q(pop_v[0]) );
  arbiter2_15 arbiter_n ( .clk(clk), .rst(rst), .request({\request[0][1] , 
        \request[0][0] }), .buffer_full_i(buffer_full_in[0]), .grant(grant_0), 
        .grant_v_o(grant_v[0]) );
  arbiter2_14 arbiter_s ( .clk(clk), .rst(rst), .request({\request[1][1] , 
        \request[1][0] }), .buffer_full_i(buffer_full_in[1]), .grant(grant_1), 
        .grant_v_o(grant_v[1]) );
  arbiter3_7 arbiter_e ( .clk(clk), .rst(rst), .request({\request[2][2] , 
        \request[2][1] , \request[2][0] }), .buffer_full_i(buffer_full_in[2]), 
        .grant(grant_2), .grant_v_o(grant_v[2]) );
  arbiter3_6 arbiter_l ( .clk(clk), .rst(rst), .request({\request[3][2] , 
        \request[3][1] , \request[3][0] }), .buffer_full_i(buffer_full_in[3]), 
        .grant({\grant_3[2] , grant_3[1:0]}), .grant_v_o(grant_v[3]) );
  dccl_35 dccl_n ( .packet_addr_y_i({\packet_addr[0][3] , \packet_addr[0][2] , 
        \packet_addr[0][1] , \packet_addr[0][0] }), .packet_addr_x_i({
        \packet_addr[0][7] , \packet_addr[0][6] , \packet_addr[0][5] , 
        \packet_addr[0][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[0]), 
        .east_req(\request[2][0] ), .south_req(\request[1][0] ), .local_req(
        \request[3][0] ) );
  dccl_34 dccl_s ( .packet_addr_y_i({\packet_addr[1][3] , \packet_addr[1][2] , 
        \packet_addr[1][1] , \packet_addr[1][0] }), .packet_addr_x_i({
        \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] , 
        \packet_addr[1][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[1]), 
        .north_req(\request[0][0] ), .east_req(\request[2][1] ), .local_req(
        \request[3][1] ) );
  dccl_33 dccl_e ( .packet_addr_y_i({\packet_addr[2][3] , \packet_addr[2][2] , 
        \packet_addr[2][1] , \packet_addr[2][0] }), .packet_addr_x_i({
        \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] , 
        \packet_addr[2][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[2]), 
        .local_req(\request[3][2] ) );
  dccl_32 dccl_l ( .packet_addr_y_i({\packet_addr[3][3] , \packet_addr[3][2] , 
        \packet_addr[3][1] , \packet_addr[3][0] }), .packet_addr_x_i({
        \packet_addr[3][7] , \packet_addr[3][6] , \packet_addr[3][5] , 
        \packet_addr[3][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[3]), 
        .north_req(\request[0][1] ), .east_req(\request[2][2] ), .south_req(
        \request[1][1] ) );
endmodule


module mux2_1_15 ( data0, data1, select0, select1, data_o );
  input [15:0] data0;
  input [15:0] data1;
  output [15:0] data_o;
  input select0, select1;
  wire   n1, n4, n5;

  AO22X1 U4 ( .IN1(data1[9]), .IN2(n5), .IN3(data0[9]), .IN4(n4), .Q(data_o[9]) );
  AO22X1 U5 ( .IN1(data1[8]), .IN2(n5), .IN3(data0[8]), .IN4(n4), .Q(data_o[8]) );
  AO22X1 U6 ( .IN1(data1[7]), .IN2(n5), .IN3(data0[7]), .IN4(n4), .Q(data_o[7]) );
  AO22X1 U7 ( .IN1(data1[6]), .IN2(n5), .IN3(data0[6]), .IN4(n4), .Q(data_o[6]) );
  AO22X1 U8 ( .IN1(data1[5]), .IN2(n5), .IN3(data0[5]), .IN4(n4), .Q(data_o[5]) );
  AO22X1 U9 ( .IN1(data1[4]), .IN2(n5), .IN3(data0[4]), .IN4(n4), .Q(data_o[4]) );
  AO22X1 U10 ( .IN1(data1[3]), .IN2(n5), .IN3(data0[3]), .IN4(n4), .Q(
        data_o[3]) );
  AO22X1 U11 ( .IN1(data1[2]), .IN2(n5), .IN3(data0[2]), .IN4(n4), .Q(
        data_o[2]) );
  AO22X1 U12 ( .IN1(data1[1]), .IN2(n5), .IN3(data0[1]), .IN4(n4), .Q(
        data_o[1]) );
  AO22X1 U13 ( .IN1(data1[15]), .IN2(n5), .IN3(data0[15]), .IN4(n4), .Q(
        data_o[15]) );
  AO22X1 U14 ( .IN1(data1[14]), .IN2(n5), .IN3(data0[14]), .IN4(n4), .Q(
        data_o[14]) );
  AO22X1 U15 ( .IN1(data1[13]), .IN2(n5), .IN3(data0[13]), .IN4(n4), .Q(
        data_o[13]) );
  AO22X1 U16 ( .IN1(data1[12]), .IN2(n5), .IN3(data0[12]), .IN4(n4), .Q(
        data_o[12]) );
  AO22X1 U17 ( .IN1(data1[11]), .IN2(n5), .IN3(data0[11]), .IN4(n4), .Q(
        data_o[11]) );
  AO22X1 U18 ( .IN1(data1[10]), .IN2(n5), .IN3(data0[10]), .IN4(n4), .Q(
        data_o[10]) );
  AO22X1 U19 ( .IN1(data1[0]), .IN2(n5), .IN3(data0[0]), .IN4(n4), .Q(
        data_o[0]) );
  INVX0 U2 ( .INP(select1), .ZN(n1) );
  AND2X1 U3 ( .IN1(select0), .IN2(n1), .Q(n4) );
  NOR2X0 U20 ( .IN1(n1), .IN2(select0), .QN(n5) );
endmodule


module mux2_1_14 ( data0, data1, select0, select1, data_o );
  input [15:0] data0;
  input [15:0] data1;
  output [15:0] data_o;
  input select0, select1;
  wire   n1, n4, n5;

  AO22X1 U4 ( .IN1(data1[9]), .IN2(n5), .IN3(data0[9]), .IN4(n4), .Q(data_o[9]) );
  AO22X1 U5 ( .IN1(data1[8]), .IN2(n5), .IN3(data0[8]), .IN4(n4), .Q(data_o[8]) );
  AO22X1 U6 ( .IN1(data1[7]), .IN2(n5), .IN3(data0[7]), .IN4(n4), .Q(data_o[7]) );
  AO22X1 U7 ( .IN1(data1[6]), .IN2(n5), .IN3(data0[6]), .IN4(n4), .Q(data_o[6]) );
  AO22X1 U8 ( .IN1(data1[5]), .IN2(n5), .IN3(data0[5]), .IN4(n4), .Q(data_o[5]) );
  AO22X1 U9 ( .IN1(data1[4]), .IN2(n5), .IN3(data0[4]), .IN4(n4), .Q(data_o[4]) );
  AO22X1 U10 ( .IN1(data1[3]), .IN2(n5), .IN3(data0[3]), .IN4(n4), .Q(
        data_o[3]) );
  AO22X1 U11 ( .IN1(data1[2]), .IN2(n5), .IN3(data0[2]), .IN4(n4), .Q(
        data_o[2]) );
  AO22X1 U12 ( .IN1(data1[1]), .IN2(n5), .IN3(data0[1]), .IN4(n4), .Q(
        data_o[1]) );
  AO22X1 U13 ( .IN1(data1[15]), .IN2(n5), .IN3(data0[15]), .IN4(n4), .Q(
        data_o[15]) );
  AO22X1 U14 ( .IN1(data1[14]), .IN2(n5), .IN3(data0[14]), .IN4(n4), .Q(
        data_o[14]) );
  AO22X1 U15 ( .IN1(data1[13]), .IN2(n5), .IN3(data0[13]), .IN4(n4), .Q(
        data_o[13]) );
  AO22X1 U16 ( .IN1(data1[12]), .IN2(n5), .IN3(data0[12]), .IN4(n4), .Q(
        data_o[12]) );
  AO22X1 U17 ( .IN1(data1[11]), .IN2(n5), .IN3(data0[11]), .IN4(n4), .Q(
        data_o[11]) );
  AO22X1 U18 ( .IN1(data1[10]), .IN2(n5), .IN3(data0[10]), .IN4(n4), .Q(
        data_o[10]) );
  AO22X1 U19 ( .IN1(data1[0]), .IN2(n5), .IN3(data0[0]), .IN4(n4), .Q(
        data_o[0]) );
  INVX0 U2 ( .INP(select1), .ZN(n1) );
  AND2X1 U3 ( .IN1(select0), .IN2(n1), .Q(n4) );
  NOR2X0 U20 ( .IN1(n1), .IN2(select0), .QN(n5) );
endmodule


module mux3_1_7 ( data0, data1, data2, select0, select1, select2, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  output [15:0] data_o;
  input select0, select1, select2;
  wire   n1, n2, n6, n7, n8;

  AO222X1 U4 ( .IN1(data1[9]), .IN2(n8), .IN3(data0[9]), .IN4(n7), .IN5(
        data2[9]), .IN6(n6), .Q(data_o[9]) );
  AO222X1 U5 ( .IN1(data1[8]), .IN2(n8), .IN3(data0[8]), .IN4(n7), .IN5(
        data2[8]), .IN6(n6), .Q(data_o[8]) );
  AO222X1 U6 ( .IN1(data1[7]), .IN2(n8), .IN3(data0[7]), .IN4(n7), .IN5(
        data2[7]), .IN6(n6), .Q(data_o[7]) );
  AO222X1 U7 ( .IN1(data1[6]), .IN2(n8), .IN3(data0[6]), .IN4(n7), .IN5(
        data2[6]), .IN6(n6), .Q(data_o[6]) );
  AO222X1 U8 ( .IN1(data1[5]), .IN2(n8), .IN3(data0[5]), .IN4(n7), .IN5(
        data2[5]), .IN6(n6), .Q(data_o[5]) );
  AO222X1 U9 ( .IN1(data1[4]), .IN2(n8), .IN3(data0[4]), .IN4(n7), .IN5(
        data2[4]), .IN6(n6), .Q(data_o[4]) );
  AO222X1 U10 ( .IN1(data1[3]), .IN2(n8), .IN3(data0[3]), .IN4(n7), .IN5(
        data2[3]), .IN6(n6), .Q(data_o[3]) );
  AO222X1 U11 ( .IN1(data1[2]), .IN2(n8), .IN3(data0[2]), .IN4(n7), .IN5(
        data2[2]), .IN6(n6), .Q(data_o[2]) );
  AO222X1 U12 ( .IN1(data1[1]), .IN2(n8), .IN3(data0[1]), .IN4(n7), .IN5(
        data2[1]), .IN6(n6), .Q(data_o[1]) );
  AO222X1 U13 ( .IN1(data1[15]), .IN2(n8), .IN3(data0[15]), .IN4(n7), .IN5(
        data2[15]), .IN6(n6), .Q(data_o[15]) );
  AO222X1 U14 ( .IN1(data1[14]), .IN2(n8), .IN3(data0[14]), .IN4(n7), .IN5(
        data2[14]), .IN6(n6), .Q(data_o[14]) );
  AO222X1 U15 ( .IN1(data1[13]), .IN2(n8), .IN3(data0[13]), .IN4(n7), .IN5(
        data2[13]), .IN6(n6), .Q(data_o[13]) );
  AO222X1 U16 ( .IN1(data1[12]), .IN2(n8), .IN3(data0[12]), .IN4(n7), .IN5(
        data2[12]), .IN6(n6), .Q(data_o[12]) );
  AO222X1 U17 ( .IN1(data1[11]), .IN2(n8), .IN3(data0[11]), .IN4(n7), .IN5(
        data2[11]), .IN6(n6), .Q(data_o[11]) );
  AO222X1 U18 ( .IN1(data1[10]), .IN2(n8), .IN3(data0[10]), .IN4(n7), .IN5(
        data2[10]), .IN6(n6), .Q(data_o[10]) );
  AO222X1 U19 ( .IN1(data1[0]), .IN2(n8), .IN3(data0[0]), .IN4(n7), .IN5(
        data2[0]), .IN6(n6), .Q(data_o[0]) );
  INVX0 U2 ( .INP(select0), .ZN(n2) );
  INVX0 U3 ( .INP(select1), .ZN(n1) );
  AND3X1 U20 ( .IN1(n2), .IN2(n1), .IN3(select2), .Q(n6) );
  NOR3X0 U21 ( .IN1(select1), .IN2(select2), .IN3(n2), .QN(n7) );
  NOR3X0 U22 ( .IN1(select0), .IN2(select2), .IN3(n1), .QN(n8) );
endmodule


module mux3_1_6 ( data0, data1, data2, select0, select1, select2, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  output [15:0] data_o;
  input select0, select1, select2;
  wire   n1, n2, n6, n7, n8;

  AO222X1 U4 ( .IN1(data1[9]), .IN2(n8), .IN3(data0[9]), .IN4(n7), .IN5(
        data2[9]), .IN6(n6), .Q(data_o[9]) );
  AO222X1 U5 ( .IN1(data1[8]), .IN2(n8), .IN3(data0[8]), .IN4(n7), .IN5(
        data2[8]), .IN6(n6), .Q(data_o[8]) );
  AO222X1 U6 ( .IN1(data1[7]), .IN2(n8), .IN3(data0[7]), .IN4(n7), .IN5(
        data2[7]), .IN6(n6), .Q(data_o[7]) );
  AO222X1 U7 ( .IN1(data1[6]), .IN2(n8), .IN3(data0[6]), .IN4(n7), .IN5(
        data2[6]), .IN6(n6), .Q(data_o[6]) );
  AO222X1 U8 ( .IN1(data1[5]), .IN2(n8), .IN3(data0[5]), .IN4(n7), .IN5(
        data2[5]), .IN6(n6), .Q(data_o[5]) );
  AO222X1 U9 ( .IN1(data1[4]), .IN2(n8), .IN3(data0[4]), .IN4(n7), .IN5(
        data2[4]), .IN6(n6), .Q(data_o[4]) );
  AO222X1 U10 ( .IN1(data1[3]), .IN2(n8), .IN3(data0[3]), .IN4(n7), .IN5(
        data2[3]), .IN6(n6), .Q(data_o[3]) );
  AO222X1 U11 ( .IN1(data1[2]), .IN2(n8), .IN3(data0[2]), .IN4(n7), .IN5(
        data2[2]), .IN6(n6), .Q(data_o[2]) );
  AO222X1 U12 ( .IN1(data1[1]), .IN2(n8), .IN3(data0[1]), .IN4(n7), .IN5(
        data2[1]), .IN6(n6), .Q(data_o[1]) );
  AO222X1 U13 ( .IN1(data1[15]), .IN2(n8), .IN3(data0[15]), .IN4(n7), .IN5(
        data2[15]), .IN6(n6), .Q(data_o[15]) );
  AO222X1 U14 ( .IN1(data1[14]), .IN2(n8), .IN3(data0[14]), .IN4(n7), .IN5(
        data2[14]), .IN6(n6), .Q(data_o[14]) );
  AO222X1 U15 ( .IN1(data1[13]), .IN2(n8), .IN3(data0[13]), .IN4(n7), .IN5(
        data2[13]), .IN6(n6), .Q(data_o[13]) );
  AO222X1 U16 ( .IN1(data1[12]), .IN2(n8), .IN3(data0[12]), .IN4(n7), .IN5(
        data2[12]), .IN6(n6), .Q(data_o[12]) );
  AO222X1 U17 ( .IN1(data1[11]), .IN2(n8), .IN3(data0[11]), .IN4(n7), .IN5(
        data2[11]), .IN6(n6), .Q(data_o[11]) );
  AO222X1 U18 ( .IN1(data1[10]), .IN2(n8), .IN3(data0[10]), .IN4(n7), .IN5(
        data2[10]), .IN6(n6), .Q(data_o[10]) );
  AO222X1 U19 ( .IN1(data1[0]), .IN2(n8), .IN3(data0[0]), .IN4(n7), .IN5(
        data2[0]), .IN6(n6), .Q(data_o[0]) );
  INVX0 U2 ( .INP(select0), .ZN(n2) );
  INVX0 U3 ( .INP(select1), .ZN(n1) );
  AND3X1 U20 ( .IN1(n2), .IN2(n1), .IN3(select2), .Q(n6) );
  NOR3X0 U21 ( .IN1(select1), .IN2(select2), .IN3(n2), .QN(n7) );
  NOR3X0 U22 ( .IN1(select0), .IN2(select2), .IN3(n1), .QN(n8) );
endmodule



    module node4_NODE_X0_NODE_Y1I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__I_node_2_node_interface__ ( 
        \clk.clk , \reset.reset , \local_node.clk , 
        \local_node.buffer_full_in , \local_node.buffer_full_out , 
        \local_node.receiving_data , \local_node.sending_data , 
        \local_node.data_in , \local_node.data_out , \node_0.clk , 
        \node_0.buffer_full_in , \node_0.buffer_full_out , 
        \node_0.receiving_data , \node_0.sending_data , \node_0.data_in , 
        \node_0.data_out , \node_1.clk , \node_1.buffer_full_in , 
        \node_1.buffer_full_out , \node_1.receiving_data , 
        \node_1.sending_data , \node_1.data_in , \node_1.data_out , 
        \node_2.clk , \node_2.buffer_full_in , \node_2.buffer_full_out , 
        \node_2.receiving_data , \node_2.sending_data , \node_2.data_in , 
        \node_2.data_out  );
  input [15:0] \local_node.data_in ;
  output [15:0] \local_node.data_out ;
  input [15:0] \node_0.data_in ;
  output [15:0] \node_0.data_out ;
  input [15:0] \node_1.data_in ;
  output [15:0] \node_1.data_out ;
  input [15:0] \node_2.data_in ;
  output [15:0] \node_2.data_out ;
  input \clk.clk , \reset.reset , \local_node.buffer_full_in ,
         \local_node.receiving_data , \node_0.buffer_full_in ,
         \node_0.receiving_data , \node_1.buffer_full_in ,
         \node_1.receiving_data , \node_2.buffer_full_in ,
         \node_2.receiving_data ;
  output \local_node.buffer_full_out , \local_node.sending_data ,
         \node_0.buffer_full_out , \node_0.sending_data ,
         \node_1.buffer_full_out , \node_1.sending_data ,
         \node_2.buffer_full_out , \node_2.sending_data ;
  inout \local_node.clk ,  \node_0.clk ,  \node_1.clk ,  \node_2.clk ;
  wire   \buffer_out[3][15] , \buffer_out[3][14] , \buffer_out[3][13] ,
         \buffer_out[3][12] , \buffer_out[3][11] , \buffer_out[3][10] ,
         \buffer_out[3][9] , \buffer_out[3][8] , \buffer_out[3][7] ,
         \buffer_out[3][6] , \buffer_out[3][5] , \buffer_out[3][4] ,
         \buffer_out[3][3] , \buffer_out[3][2] , \buffer_out[3][1] ,
         \buffer_out[3][0] , \buffer_out[2][15] , \buffer_out[2][14] ,
         \buffer_out[2][13] , \buffer_out[2][12] , \buffer_out[2][11] ,
         \buffer_out[2][10] , \buffer_out[2][9] , \buffer_out[2][8] ,
         \buffer_out[2][7] , \buffer_out[2][6] , \buffer_out[2][5] ,
         \buffer_out[2][4] , \buffer_out[2][3] , \buffer_out[2][2] ,
         \buffer_out[2][1] , \buffer_out[2][0] , \buffer_out[1][15] ,
         \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] ,
         \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] ,
         \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] ,
         \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] ,
         \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] ,
         \buffer_out[0][15] , \buffer_out[0][14] , \buffer_out[0][13] ,
         \buffer_out[0][12] , \buffer_out[0][11] , \buffer_out[0][10] ,
         \buffer_out[0][9] , \buffer_out[0][8] , \buffer_out[0][7] ,
         \buffer_out[0][6] , \buffer_out[0][5] , \buffer_out[0][4] ,
         \buffer_out[0][3] , \buffer_out[0][2] , \buffer_out[0][1] ,
         \buffer_out[0][0] , \next_buffer_out[3][15] ,
         \next_buffer_out[3][14] , \next_buffer_out[3][13] ,
         \next_buffer_out[3][12] , \next_buffer_out[3][11] ,
         \next_buffer_out[3][10] , \next_buffer_out[3][9] ,
         \next_buffer_out[3][8] , \next_buffer_out[3][7] ,
         \next_buffer_out[3][6] , \next_buffer_out[3][5] ,
         \next_buffer_out[3][4] , \next_buffer_out[3][3] ,
         \next_buffer_out[3][2] , \next_buffer_out[3][1] ,
         \next_buffer_out[3][0] , \next_buffer_out[2][15] ,
         \next_buffer_out[2][14] , \next_buffer_out[2][13] ,
         \next_buffer_out[2][12] , \next_buffer_out[2][11] ,
         \next_buffer_out[2][10] , \next_buffer_out[2][9] ,
         \next_buffer_out[2][8] , \next_buffer_out[2][7] ,
         \next_buffer_out[2][6] , \next_buffer_out[2][5] ,
         \next_buffer_out[2][4] , \next_buffer_out[2][3] ,
         \next_buffer_out[2][2] , \next_buffer_out[2][1] ,
         \next_buffer_out[2][0] , \next_buffer_out[1][15] ,
         \next_buffer_out[1][14] , \next_buffer_out[1][13] ,
         \next_buffer_out[1][12] , \next_buffer_out[1][11] ,
         \next_buffer_out[1][10] , \next_buffer_out[1][9] ,
         \next_buffer_out[1][8] , \next_buffer_out[1][7] ,
         \next_buffer_out[1][6] , \next_buffer_out[1][5] ,
         \next_buffer_out[1][4] , \next_buffer_out[1][3] ,
         \next_buffer_out[1][2] , \next_buffer_out[1][1] ,
         \next_buffer_out[1][0] , \next_buffer_out[0][15] ,
         \next_buffer_out[0][14] , \next_buffer_out[0][13] ,
         \next_buffer_out[0][12] , \next_buffer_out[0][11] ,
         \next_buffer_out[0][10] , \next_buffer_out[0][9] ,
         \next_buffer_out[0][8] , \next_buffer_out[0][7] ,
         \next_buffer_out[0][6] , \next_buffer_out[0][5] ,
         \next_buffer_out[0][4] , \next_buffer_out[0][3] ,
         \next_buffer_out[0][2] , \next_buffer_out[0][1] ,
         \next_buffer_out[0][0] ;
  wire   [3:0] buffer_full_in;
  wire   [3:0] receiving_data;
  wire   [3:0] pop_v;
  wire   [3:0] data_valid;
  wire   [3:0] next_data_valid;
  wire   [1:0] grant_0;
  wire   [1:0] grant_1;
  wire   [2:0] grant_2;
  wire   [2:0] grant_3;
  tri   \local_node.buffer_full_in ;
  tri   \local_node.buffer_full_out ;
  tri   \local_node.receiving_data ;
  tri   \local_node.sending_data ;
  tri   [15:0] \local_node.data_in ;
  tri   [15:0] \local_node.data_out ;

  converter_out_I_n_node_interface_dut_ c3 ( .\n.buffer_full_in (
        \local_node.buffer_full_in ), .\n.receiving_data (
        \local_node.receiving_data ), .\n.data_in (\local_node.data_in ), 
        .\n.buffer_full_out (\local_node.buffer_full_out ), .\n.sending_data (
        \local_node.sending_data ), .\n.data_out (\local_node.data_out ), 
        .buffer_full_in(1'b0), .receiving_data(1'b0), .data_in({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  fifo_kev_35 \genblk1[0].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[0]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[0]), .data_out({\buffer_out[0][15] , 
        \buffer_out[0][14] , \buffer_out[0][13] , \buffer_out[0][12] , 
        \buffer_out[0][11] , \buffer_out[0][10] , \buffer_out[0][9] , 
        \buffer_out[0][8] , \buffer_out[0][7] , \buffer_out[0][6] , 
        \buffer_out[0][5] , \buffer_out[0][4] , \buffer_out[0][3] , 
        \buffer_out[0][2] , \buffer_out[0][1] , \buffer_out[0][0] }), 
        .next_data_out({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] , 
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .next_data_valid(
        next_data_valid[0]) );
  address_counter_35 \genblk1[0].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] }), 
        .buffer_data_valid(next_data_valid[0]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .buffer_pop(
        pop_v[0]), .receiving_data(1'b0) );
  fifo_kev_34 \genblk1[1].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[1]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[1]), .data_out({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), 
        .next_data_out({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] , 
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .next_data_valid(
        next_data_valid[1]) );
  address_counter_34 \genblk1[1].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] }), 
        .buffer_data_valid(next_data_valid[1]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .buffer_pop(
        pop_v[1]), .receiving_data(1'b0) );
  fifo_kev_33 \genblk1[2].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[2]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[2]), .data_out({\buffer_out[2][15] , 
        \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] , 
        \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] , 
        \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] , 
        \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] , 
        \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] }), 
        .next_data_out({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] , 
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .next_data_valid(
        next_data_valid[2]) );
  address_counter_33 \genblk1[2].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] }), 
        .buffer_data_valid(next_data_valid[2]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .buffer_pop(
        pop_v[2]), .receiving_data(1'b0) );
  fifo_kev_32 \genblk1[3].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[3]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[3]), .data_out({\buffer_out[3][15] , 
        \buffer_out[3][14] , \buffer_out[3][13] , \buffer_out[3][12] , 
        \buffer_out[3][11] , \buffer_out[3][10] , \buffer_out[3][9] , 
        \buffer_out[3][8] , \buffer_out[3][7] , \buffer_out[3][6] , 
        \buffer_out[3][5] , \buffer_out[3][4] , \buffer_out[3][3] , 
        \buffer_out[3][2] , \buffer_out[3][1] , \buffer_out[3][0] }), 
        .next_data_out({\next_buffer_out[3][15] , \next_buffer_out[3][14] , 
        \next_buffer_out[3][13] , \next_buffer_out[3][12] , 
        \next_buffer_out[3][11] , \next_buffer_out[3][10] , 
        \next_buffer_out[3][9] , \next_buffer_out[3][8] , 
        \next_buffer_out[3][7] , \next_buffer_out[3][6] , 
        \next_buffer_out[3][5] , \next_buffer_out[3][4] , 
        \next_buffer_out[3][3] , \next_buffer_out[3][2] , 
        \next_buffer_out[3][1] , \next_buffer_out[3][0] }), .next_data_valid(
        next_data_valid[3]) );
  address_counter_32 \genblk1[3].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[3][15] , \next_buffer_out[3][14] , 
        \next_buffer_out[3][13] , \next_buffer_out[3][12] , 
        \next_buffer_out[3][11] , \next_buffer_out[3][10] , 
        \next_buffer_out[3][9] , \next_buffer_out[3][8] }), 
        .buffer_data_valid(next_data_valid[3]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[3][7] , \next_buffer_out[3][6] , 
        \next_buffer_out[3][5] , \next_buffer_out[3][4] , 
        \next_buffer_out[3][3] , \next_buffer_out[3][2] , 
        \next_buffer_out[3][1] , \next_buffer_out[3][0] }), .buffer_pop(
        pop_v[3]), .receiving_data(1'b0) );
  converter_in_I_n_node_interface_dut__13 \genblk2.c0  ( .\n.buffer_full_in (
        \node_0.buffer_full_in ), .\n.receiving_data (\node_0.receiving_data ), 
        .\n.data_in (\node_0.data_in ), .\n.buffer_full_out (
        \node_0.buffer_full_out ), .\n.sending_data (\node_0.sending_data ), 
        .\n.data_out (\node_0.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_out_I_n_node_interface_dut_ \genblk2.c1  ( .\n.buffer_full_in (
        \node_1.buffer_full_in ), .\n.receiving_data (\node_1.receiving_data ), 
        .\n.data_in (\node_1.data_in ), .\n.buffer_full_out (
        \node_1.buffer_full_out ), .\n.sending_data (\node_1.sending_data ), 
        .\n.data_out (\node_1.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_in_I_n_node_interface_dut__12 \genblk2.c2  ( .\n.buffer_full_in (
        \node_2.buffer_full_in ), .\n.receiving_data (\node_2.receiving_data ), 
        .\n.data_in (\node_2.data_in ), .\n.buffer_full_out (
        \node_2.buffer_full_out ), .\n.sending_data (\node_2.sending_data ), 
        .\n.data_out (\node_2.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  controller4_edge_w_1 \genblk2.w  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .packet_addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .local_addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), 
        .packet_valid(data_valid), .buffer_full_in({1'b0, 1'b0, 1'b0, 1'b0}), 
        .grant_0(grant_0), .grant_1(grant_1), .grant_2(grant_2), .grant_3(
        grant_3), .pop_v(pop_v) );
  mux2_1_15 \genblk2.mux_n  ( .data0({\buffer_out[1][15] , \buffer_out[1][14] , 
        \buffer_out[1][13] , \buffer_out[1][12] , \buffer_out[1][11] , 
        \buffer_out[1][10] , \buffer_out[1][9] , \buffer_out[1][8] , 
        \buffer_out[1][7] , \buffer_out[1][6] , \buffer_out[1][5] , 
        \buffer_out[1][4] , \buffer_out[1][3] , \buffer_out[1][2] , 
        \buffer_out[1][1] , \buffer_out[1][0] }), .data1({\buffer_out[3][15] , 
        \buffer_out[3][14] , \buffer_out[3][13] , \buffer_out[3][12] , 
        \buffer_out[3][11] , \buffer_out[3][10] , \buffer_out[3][9] , 
        \buffer_out[3][8] , \buffer_out[3][7] , \buffer_out[3][6] , 
        \buffer_out[3][5] , \buffer_out[3][4] , \buffer_out[3][3] , 
        \buffer_out[3][2] , \buffer_out[3][1] , \buffer_out[3][0] }), 
        .select0(grant_0[0]), .select1(grant_0[1]) );
  mux2_1_14 \genblk2.mux_s  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[3][15] , 
        \buffer_out[3][14] , \buffer_out[3][13] , \buffer_out[3][12] , 
        \buffer_out[3][11] , \buffer_out[3][10] , \buffer_out[3][9] , 
        \buffer_out[3][8] , \buffer_out[3][7] , \buffer_out[3][6] , 
        \buffer_out[3][5] , \buffer_out[3][4] , \buffer_out[3][3] , 
        \buffer_out[3][2] , \buffer_out[3][1] , \buffer_out[3][0] }), 
        .select0(grant_1[0]), .select1(grant_1[1]) );
  mux3_1_7 \genblk2.mux_e  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[3][15] , \buffer_out[3][14] , \buffer_out[3][13] , 
        \buffer_out[3][12] , \buffer_out[3][11] , \buffer_out[3][10] , 
        \buffer_out[3][9] , \buffer_out[3][8] , \buffer_out[3][7] , 
        \buffer_out[3][6] , \buffer_out[3][5] , \buffer_out[3][4] , 
        \buffer_out[3][3] , \buffer_out[3][2] , \buffer_out[3][1] , 
        \buffer_out[3][0] }), .select0(grant_2[0]), .select1(grant_2[1]), 
        .select2(grant_2[2]) );
  mux3_1_6 \genblk2.mux_l  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[2][15] , \buffer_out[2][14] , \buffer_out[2][13] , 
        \buffer_out[2][12] , \buffer_out[2][11] , \buffer_out[2][10] , 
        \buffer_out[2][9] , \buffer_out[2][8] , \buffer_out[2][7] , 
        \buffer_out[2][6] , \buffer_out[2][5] , \buffer_out[2][4] , 
        \buffer_out[2][3] , \buffer_out[2][2] , \buffer_out[2][1] , 
        \buffer_out[2][0] }), .select0(grant_3[0]), .select1(grant_3[1]), 
        .select2(grant_3[2]) );
endmodule


module fifo_kev_31 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_63 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_31 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_63 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_62 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_31 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_62 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_31_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_31 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_31 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_31 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_31_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_30 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_61 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_30 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_61 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_60 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_30 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_60 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_30_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_30 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_30 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_30 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_30_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_29 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_59 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_29 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_59 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_58 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_29 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_58 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_29_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_29 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_29 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_29 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_29_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_28 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_57 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_28 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_57 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_56 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_28 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_56 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_28_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_28 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_28 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_28 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_28_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module converter_in_I_n_node_interface_dut__11 ( \n.buffer_full_in , 
        \n.receiving_data , \n.data_in , \n.buffer_full_out , \n.sending_data , 
        \n.data_out , buffer_full_out, sending_data, data_out, buffer_full_in, 
        receiving_data, data_in );
  input [15:0] \n.data_in ;
  output [15:0] \n.data_out ;
  output [15:0] data_out;
  input [15:0] data_in;
  input \n.buffer_full_in , \n.receiving_data , buffer_full_in, receiving_data;
  output \n.buffer_full_out , \n.sending_data , buffer_full_out, sending_data;
  wire   \n.buffer_full_in , \n.receiving_data , buffer_full_in,
         receiving_data;
  assign buffer_full_out = \n.buffer_full_in ;
  assign sending_data = \n.receiving_data ;
  assign data_out[15] = \n.data_in  [15];
  assign data_out[14] = \n.data_in  [14];
  assign data_out[13] = \n.data_in  [13];
  assign data_out[12] = \n.data_in  [12];
  assign data_out[11] = \n.data_in  [11];
  assign data_out[10] = \n.data_in  [10];
  assign data_out[9] = \n.data_in  [9];
  assign data_out[8] = \n.data_in  [8];
  assign data_out[7] = \n.data_in  [7];
  assign data_out[6] = \n.data_in  [6];
  assign data_out[5] = \n.data_in  [5];
  assign data_out[4] = \n.data_in  [4];
  assign data_out[3] = \n.data_in  [3];
  assign data_out[2] = \n.data_in  [2];
  assign data_out[1] = \n.data_in  [1];
  assign data_out[0] = \n.data_in  [0];
  assign \n.buffer_full_out  = buffer_full_in;
  assign \n.sending_data  = receiving_data;
  assign \n.data_out  [15] = data_in[15];
  assign \n.data_out  [14] = data_in[14];
  assign \n.data_out  [13] = data_in[13];
  assign \n.data_out  [12] = data_in[12];
  assign \n.data_out  [11] = data_in[11];
  assign \n.data_out  [10] = data_in[10];
  assign \n.data_out  [9] = data_in[9];
  assign \n.data_out  [8] = data_in[8];
  assign \n.data_out  [7] = data_in[7];
  assign \n.data_out  [6] = data_in[6];
  assign \n.data_out  [5] = data_in[5];
  assign \n.data_out  [4] = data_in[4];
  assign \n.data_out  [3] = data_in[3];
  assign \n.data_out  [2] = data_in[2];
  assign \n.data_out  [1] = data_in[1];
  assign \n.data_out  [0] = data_in[0];

endmodule


module converter_in_I_n_node_interface_dut__10 ( \n.buffer_full_in , 
        \n.receiving_data , \n.data_in , \n.buffer_full_out , \n.sending_data , 
        \n.data_out , buffer_full_out, sending_data, data_out, buffer_full_in, 
        receiving_data, data_in );
  input [15:0] \n.data_in ;
  output [15:0] \n.data_out ;
  output [15:0] data_out;
  input [15:0] data_in;
  input \n.buffer_full_in , \n.receiving_data , buffer_full_in, receiving_data;
  output \n.buffer_full_out , \n.sending_data , buffer_full_out, sending_data;
  wire   \n.buffer_full_in , \n.receiving_data , buffer_full_in,
         receiving_data;
  assign buffer_full_out = \n.buffer_full_in ;
  assign sending_data = \n.receiving_data ;
  assign data_out[15] = \n.data_in  [15];
  assign data_out[14] = \n.data_in  [14];
  assign data_out[13] = \n.data_in  [13];
  assign data_out[12] = \n.data_in  [12];
  assign data_out[11] = \n.data_in  [11];
  assign data_out[10] = \n.data_in  [10];
  assign data_out[9] = \n.data_in  [9];
  assign data_out[8] = \n.data_in  [8];
  assign data_out[7] = \n.data_in  [7];
  assign data_out[6] = \n.data_in  [6];
  assign data_out[5] = \n.data_in  [5];
  assign data_out[4] = \n.data_in  [4];
  assign data_out[3] = \n.data_in  [3];
  assign data_out[2] = \n.data_in  [2];
  assign data_out[1] = \n.data_in  [1];
  assign data_out[0] = \n.data_in  [0];
  assign \n.buffer_full_out  = buffer_full_in;
  assign \n.sending_data  = receiving_data;
  assign \n.data_out  [15] = data_in[15];
  assign \n.data_out  [14] = data_in[14];
  assign \n.data_out  [13] = data_in[13];
  assign \n.data_out  [12] = data_in[12];
  assign \n.data_out  [11] = data_in[11];
  assign \n.data_out  [10] = data_in[10];
  assign \n.data_out  [9] = data_in[9];
  assign \n.data_out  [8] = data_in[8];
  assign \n.data_out  [7] = data_in[7];
  assign \n.data_out  [6] = data_in[6];
  assign \n.data_out  [5] = data_in[5];
  assign \n.data_out  [4] = data_in[4];
  assign \n.data_out  [3] = data_in[3];
  assign \n.data_out  [2] = data_in[2];
  assign \n.data_out  [1] = data_in[1];
  assign \n.data_out  [0] = data_in[0];

endmodule


module flipflop_BITS2_13 ( clk, data_i, data_o );
  input [1:0] data_i;
  output [1:0] data_o;
  input clk;


  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS2_13 ( clk, enable_i, reset, data_i, data_o );
  input [1:0] data_i;
  input [1:0] data_o;
  input clk, enable_i, reset;
  wire   n10, n11, n1, n5, n7, n8, n9;
  wire   [1:0] write_data;

  AOI22X1 U5 ( .IN1(enable_i), .IN2(data_i[1]), .IN3(n10), .IN4(n1), .QN(n9)
         );
  AOI22X1 U6 ( .IN1(data_i[0]), .IN2(enable_i), .IN3(n11), .IN4(n1), .QN(n8)
         );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n9), .QN(write_data[1]) );
  NOR2X0 U4 ( .IN1(reset), .IN2(n8), .QN(write_data[0]) );
  AND2X1 U7 ( .IN1(data_o[1]), .IN2(n7), .Q(n10) );
  AND2X1 U8 ( .IN1(data_o[0]), .IN2(n5), .Q(n11) );
  flipflop_BITS2_13 FF ( .clk(clk), .data_i(write_data), .data_o({n7, n5}) );
endmodule


module flipflop_BITS1_49 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_49 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_49 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter2_13 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [1:0] request;
  output [1:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   tail_en, n1, n2;
  wire   [1:0] req_i;
  wire   [1:0] req_o;

  AND3X1 U10 ( .IN1(request[1]), .IN2(n1), .IN3(n2), .Q(grant[1]) );
  AND3X1 U11 ( .IN1(request[0]), .IN2(n2), .IN3(request[1]), .Q(tail_en) );
  INVX0 U6 ( .INP(request[0]), .ZN(n1) );
  NOR2X0 U7 ( .IN1(buffer_full_i), .IN2(n1), .QN(grant[0]) );
  INVX0 U8 ( .INP(buffer_full_i), .ZN(n2) );
  OA21X1 U9 ( .IN1(request[1]), .IN2(request[0]), .IN3(n2), .Q(grant_v_o) );
  register_BITS2_13 req_record ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i({1'b1, 1'b0}), .data_o({1'b0, 1'b0}) );
  register_BITS1_49 tail ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i(1'b1), .data_o(1'b0) );
endmodule


module flipflop_BITS2_12 ( clk, data_i, data_o );
  input [1:0] data_i;
  output [1:0] data_o;
  input clk;


  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS2_12 ( clk, enable_i, reset, data_i, data_o );
  input [1:0] data_i;
  input [1:0] data_o;
  input clk, enable_i, reset;
  wire   n10, n11, n1, n5, n7, n8, n9;
  wire   [1:0] write_data;

  AOI22X1 U5 ( .IN1(enable_i), .IN2(data_i[1]), .IN3(n10), .IN4(n1), .QN(n9)
         );
  AOI22X1 U6 ( .IN1(data_i[0]), .IN2(enable_i), .IN3(n11), .IN4(n1), .QN(n8)
         );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n9), .QN(write_data[1]) );
  NOR2X0 U4 ( .IN1(reset), .IN2(n8), .QN(write_data[0]) );
  AND2X1 U7 ( .IN1(data_o[1]), .IN2(n7), .Q(n10) );
  AND2X1 U8 ( .IN1(data_o[0]), .IN2(n5), .Q(n11) );
  flipflop_BITS2_12 FF ( .clk(clk), .data_i(write_data), .data_o({n7, n5}) );
endmodule


module flipflop_BITS1_48 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_48 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_48 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter2_12 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [1:0] request;
  output [1:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   tail_en, n1, n2;
  wire   [1:0] req_i;
  wire   [1:0] req_o;

  AND3X1 U10 ( .IN1(request[1]), .IN2(n1), .IN3(n2), .Q(grant[1]) );
  AND3X1 U11 ( .IN1(request[0]), .IN2(n2), .IN3(request[1]), .Q(tail_en) );
  INVX0 U6 ( .INP(request[0]), .ZN(n1) );
  NOR2X0 U7 ( .IN1(buffer_full_i), .IN2(n1), .QN(grant[0]) );
  INVX0 U8 ( .INP(buffer_full_i), .ZN(n2) );
  OA21X1 U9 ( .IN1(request[1]), .IN2(request[0]), .IN3(n2), .Q(grant_v_o) );
  register_BITS2_12 req_record ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i({1'b1, 1'b0}), .data_o({1'b0, 1'b0}) );
  register_BITS1_48 tail ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i(1'b1), .data_o(1'b0) );
endmodule


module flipflop_BITS3_11 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_11 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_11 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS3_10 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_10 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_10 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS1_47 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_47 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_47 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_46 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_46 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_46 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter3_5 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [2:0] request;
  output [2:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[1][2] , \req_i[1][1] , \req_i[1][0] , \req_i[0][2] ,
         \req_i[0][1] , tail_en, N99, N100, N101, N110, N111, N118, N119, N120,
         N121, n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [1:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N99 = request[0];
  assign N100 = request[1];
  assign N101 = request[2];

  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(N111), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(N110), .Q(\req_i[0][1] ) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N121), .D(tail_en), .Q(req_en[0]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N120), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N119), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N118), .Q(grant[0]) );
  AND2X1 U20 ( .IN1(n8), .IN2(N101), .Q(n7) );
  OR3X1 U21 ( .IN1(n3), .IN2(N111), .IN3(n6), .Q(N121) );
  NOR3X0 U22 ( .IN1(N99), .IN2(N100), .IN3(n6), .QN(N120) );
  NOR3X0 U23 ( .IN1(n2), .IN2(N99), .IN3(n6), .QN(N119) );
  NAND3X0 U24 ( .IN1(n2), .IN2(n3), .IN3(n1), .QN(n5) );
  AO22X1 U25 ( .IN1(N100), .IN2(N101), .IN3(N99), .IN4(N101), .Q(N111) );
  INVX0 U10 ( .INP(N101), .ZN(n3) );
  NAND2X1 U11 ( .IN1(n5), .IN2(n4), .QN(n6) );
  INVX0 U12 ( .INP(N99), .ZN(n1) );
  INVX0 U13 ( .INP(N100), .ZN(n2) );
  INVX0 U14 ( .INP(buffer_full_i), .ZN(n4) );
  NAND2X1 U15 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NOR2X0 U16 ( .IN1(n1), .IN2(n6), .QN(N118) );
  NOR2X0 U17 ( .IN1(n1), .IN2(n2), .QN(N110) );
  OA21X1 U18 ( .IN1(N110), .IN2(n7), .IN3(n4), .Q(tail_en) );
  OA21X1 U19 ( .IN1(N101), .IN2(n8), .IN3(n4), .Q(grant_v_o) );
  register_BITS3_11 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][2] , \req_i[0][1] , 1'b0}), .data_o({
        1'b0, 1'b0, 1'b0}) );
  register_BITS3_10 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][2] , \req_i[1][1] , \req_i[1][0] }), 
        .data_o({1'b0, 1'b0, 1'b0}) );
  register_BITS1_47 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b1), .data_o(1'b0) );
  register_BITS1_46 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module flipflop_BITS3_9 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_9 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_9 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS3_8 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_8 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_8 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS1_45 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_45 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_45 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_44 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_44 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_44 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter3_4 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [2:0] request;
  output [2:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[1][2] , \req_i[1][1] , \req_i[1][0] , \req_i[0][2] ,
         \req_i[0][1] , tail_en, N99, N100, N101, N110, N111, N118, N119, N120,
         N121, n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [1:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N99 = request[0];
  assign N100 = request[1];
  assign N101 = request[2];

  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(N111), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(N110), .Q(\req_i[0][1] ) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N121), .D(tail_en), .Q(req_en[0]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N120), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N119), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N118), .Q(grant[0]) );
  AND2X1 U20 ( .IN1(n8), .IN2(N101), .Q(n7) );
  OR3X1 U21 ( .IN1(n3), .IN2(N111), .IN3(n6), .Q(N121) );
  NOR3X0 U22 ( .IN1(N99), .IN2(N100), .IN3(n6), .QN(N120) );
  NOR3X0 U23 ( .IN1(n2), .IN2(N99), .IN3(n6), .QN(N119) );
  NAND3X0 U24 ( .IN1(n2), .IN2(n3), .IN3(n1), .QN(n5) );
  AO22X1 U25 ( .IN1(N100), .IN2(N101), .IN3(N99), .IN4(N101), .Q(N111) );
  INVX0 U10 ( .INP(N101), .ZN(n3) );
  NAND2X1 U11 ( .IN1(n5), .IN2(n4), .QN(n6) );
  INVX0 U12 ( .INP(N99), .ZN(n1) );
  INVX0 U13 ( .INP(N100), .ZN(n2) );
  INVX0 U14 ( .INP(buffer_full_i), .ZN(n4) );
  NAND2X1 U15 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NOR2X0 U16 ( .IN1(n1), .IN2(n6), .QN(N118) );
  NOR2X0 U17 ( .IN1(n1), .IN2(n2), .QN(N110) );
  OA21X1 U18 ( .IN1(N110), .IN2(n7), .IN3(n4), .Q(tail_en) );
  OA21X1 U19 ( .IN1(N101), .IN2(n8), .IN3(n4), .Q(grant_v_o) );
  register_BITS3_9 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][2] , \req_i[0][1] , 1'b0}), .data_o({
        1'b0, 1'b0, 1'b0}) );
  register_BITS3_8 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][2] , \req_i[1][1] , \req_i[1][0] }), 
        .data_o({1'b0, 1'b0, 1'b0}) );
  register_BITS1_45 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b1), .data_o(1'b0) );
  register_BITS1_44 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module dccl_31 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_30 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_29 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_28 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module controller4_edge_w_0 ( clk, rst, .packet_addr({\packet_addr[3][7] , 
        \packet_addr[3][6] , \packet_addr[3][5] , \packet_addr[3][4] , 
        \packet_addr[3][3] , \packet_addr[3][2] , \packet_addr[3][1] , 
        \packet_addr[3][0] , \packet_addr[2][7] , \packet_addr[2][6] , 
        \packet_addr[2][5] , \packet_addr[2][4] , \packet_addr[2][3] , 
        \packet_addr[2][2] , \packet_addr[2][1] , \packet_addr[2][0] , 
        \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] , 
        \packet_addr[1][4] , \packet_addr[1][3] , \packet_addr[1][2] , 
        \packet_addr[1][1] , \packet_addr[1][0] , \packet_addr[0][7] , 
        \packet_addr[0][6] , \packet_addr[0][5] , \packet_addr[0][4] , 
        \packet_addr[0][3] , \packet_addr[0][2] , \packet_addr[0][1] , 
        \packet_addr[0][0] }), local_addr, packet_valid, buffer_full_in, 
        grant_0, grant_1, grant_2, grant_3, grant_v, pop_v );
  input [7:0] local_addr;
  input [3:0] packet_valid;
  input [3:0] buffer_full_in;
  output [1:0] grant_0;
  output [1:0] grant_1;
  output [2:0] grant_2;
  output [2:0] grant_3;
  output [3:0] grant_v;
  output [3:0] pop_v;
  input clk, rst, \packet_addr[3][7] , \packet_addr[3][6] ,
         \packet_addr[3][5] , \packet_addr[3][4] , \packet_addr[3][3] ,
         \packet_addr[3][2] , \packet_addr[3][1] , \packet_addr[3][0] ,
         \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] ,
         \packet_addr[2][4] , \packet_addr[2][3] , \packet_addr[2][2] ,
         \packet_addr[2][1] , \packet_addr[2][0] , \packet_addr[1][7] ,
         \packet_addr[1][6] , \packet_addr[1][5] , \packet_addr[1][4] ,
         \packet_addr[1][3] , \packet_addr[1][2] , \packet_addr[1][1] ,
         \packet_addr[1][0] , \packet_addr[0][7] , \packet_addr[0][6] ,
         \packet_addr[0][5] , \packet_addr[0][4] , \packet_addr[0][3] ,
         \packet_addr[0][2] , \packet_addr[0][1] , \packet_addr[0][0] ;
  wire   \grant_3[2] , \request[3][2] , \request[3][1] , \request[3][0] ,
         \request[2][2] , \request[2][1] , \request[2][0] , \request[1][1] ,
         \request[1][0] , \request[0][1] , \request[0][0] ;
  assign pop_v[2] = \grant_3[2] ;
  assign grant_3[2] = \grant_3[2] ;

  OR3X1 U1 ( .IN1(grant_2[2]), .IN2(grant_1[1]), .IN3(grant_0[1]), .Q(pop_v[3]) );
  OR3X1 U2 ( .IN1(grant_3[1]), .IN2(grant_2[1]), .IN3(grant_0[0]), .Q(pop_v[1]) );
  OR3X1 U3 ( .IN1(grant_3[0]), .IN2(grant_2[0]), .IN3(grant_1[0]), .Q(pop_v[0]) );
  arbiter2_13 arbiter_n ( .clk(clk), .rst(rst), .request({\request[0][1] , 
        \request[0][0] }), .buffer_full_i(buffer_full_in[0]), .grant(grant_0), 
        .grant_v_o(grant_v[0]) );
  arbiter2_12 arbiter_s ( .clk(clk), .rst(rst), .request({\request[1][1] , 
        \request[1][0] }), .buffer_full_i(buffer_full_in[1]), .grant(grant_1), 
        .grant_v_o(grant_v[1]) );
  arbiter3_5 arbiter_e ( .clk(clk), .rst(rst), .request({\request[2][2] , 
        \request[2][1] , \request[2][0] }), .buffer_full_i(buffer_full_in[2]), 
        .grant(grant_2), .grant_v_o(grant_v[2]) );
  arbiter3_4 arbiter_l ( .clk(clk), .rst(rst), .request({\request[3][2] , 
        \request[3][1] , \request[3][0] }), .buffer_full_i(buffer_full_in[3]), 
        .grant({\grant_3[2] , grant_3[1:0]}), .grant_v_o(grant_v[3]) );
  dccl_31 dccl_n ( .packet_addr_y_i({\packet_addr[0][3] , \packet_addr[0][2] , 
        \packet_addr[0][1] , \packet_addr[0][0] }), .packet_addr_x_i({
        \packet_addr[0][7] , \packet_addr[0][6] , \packet_addr[0][5] , 
        \packet_addr[0][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[0]), 
        .east_req(\request[2][0] ), .south_req(\request[1][0] ), .local_req(
        \request[3][0] ) );
  dccl_30 dccl_s ( .packet_addr_y_i({\packet_addr[1][3] , \packet_addr[1][2] , 
        \packet_addr[1][1] , \packet_addr[1][0] }), .packet_addr_x_i({
        \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] , 
        \packet_addr[1][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[1]), 
        .north_req(\request[0][0] ), .east_req(\request[2][1] ), .local_req(
        \request[3][1] ) );
  dccl_29 dccl_e ( .packet_addr_y_i({\packet_addr[2][3] , \packet_addr[2][2] , 
        \packet_addr[2][1] , \packet_addr[2][0] }), .packet_addr_x_i({
        \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] , 
        \packet_addr[2][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[2]), 
        .local_req(\request[3][2] ) );
  dccl_28 dccl_l ( .packet_addr_y_i({\packet_addr[3][3] , \packet_addr[3][2] , 
        \packet_addr[3][1] , \packet_addr[3][0] }), .packet_addr_x_i({
        \packet_addr[3][7] , \packet_addr[3][6] , \packet_addr[3][5] , 
        \packet_addr[3][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[3]), 
        .north_req(\request[0][1] ), .east_req(\request[2][2] ), .south_req(
        \request[1][1] ) );
endmodule


module mux2_1_13 ( data0, data1, select0, select1, data_o );
  input [15:0] data0;
  input [15:0] data1;
  output [15:0] data_o;
  input select0, select1;
  wire   n1, n4, n5;

  AO22X1 U4 ( .IN1(data1[9]), .IN2(n5), .IN3(data0[9]), .IN4(n4), .Q(data_o[9]) );
  AO22X1 U5 ( .IN1(data1[8]), .IN2(n5), .IN3(data0[8]), .IN4(n4), .Q(data_o[8]) );
  AO22X1 U6 ( .IN1(data1[7]), .IN2(n5), .IN3(data0[7]), .IN4(n4), .Q(data_o[7]) );
  AO22X1 U7 ( .IN1(data1[6]), .IN2(n5), .IN3(data0[6]), .IN4(n4), .Q(data_o[6]) );
  AO22X1 U8 ( .IN1(data1[5]), .IN2(n5), .IN3(data0[5]), .IN4(n4), .Q(data_o[5]) );
  AO22X1 U9 ( .IN1(data1[4]), .IN2(n5), .IN3(data0[4]), .IN4(n4), .Q(data_o[4]) );
  AO22X1 U10 ( .IN1(data1[3]), .IN2(n5), .IN3(data0[3]), .IN4(n4), .Q(
        data_o[3]) );
  AO22X1 U11 ( .IN1(data1[2]), .IN2(n5), .IN3(data0[2]), .IN4(n4), .Q(
        data_o[2]) );
  AO22X1 U12 ( .IN1(data1[1]), .IN2(n5), .IN3(data0[1]), .IN4(n4), .Q(
        data_o[1]) );
  AO22X1 U13 ( .IN1(data1[15]), .IN2(n5), .IN3(data0[15]), .IN4(n4), .Q(
        data_o[15]) );
  AO22X1 U14 ( .IN1(data1[14]), .IN2(n5), .IN3(data0[14]), .IN4(n4), .Q(
        data_o[14]) );
  AO22X1 U15 ( .IN1(data1[13]), .IN2(n5), .IN3(data0[13]), .IN4(n4), .Q(
        data_o[13]) );
  AO22X1 U16 ( .IN1(data1[12]), .IN2(n5), .IN3(data0[12]), .IN4(n4), .Q(
        data_o[12]) );
  AO22X1 U17 ( .IN1(data1[11]), .IN2(n5), .IN3(data0[11]), .IN4(n4), .Q(
        data_o[11]) );
  AO22X1 U18 ( .IN1(data1[10]), .IN2(n5), .IN3(data0[10]), .IN4(n4), .Q(
        data_o[10]) );
  AO22X1 U19 ( .IN1(data1[0]), .IN2(n5), .IN3(data0[0]), .IN4(n4), .Q(
        data_o[0]) );
  INVX0 U2 ( .INP(select1), .ZN(n1) );
  AND2X1 U3 ( .IN1(select0), .IN2(n1), .Q(n4) );
  NOR2X0 U20 ( .IN1(n1), .IN2(select0), .QN(n5) );
endmodule


module mux2_1_12 ( data0, data1, select0, select1, data_o );
  input [15:0] data0;
  input [15:0] data1;
  output [15:0] data_o;
  input select0, select1;
  wire   n1, n4, n5;

  AO22X1 U4 ( .IN1(data1[9]), .IN2(n5), .IN3(data0[9]), .IN4(n4), .Q(data_o[9]) );
  AO22X1 U5 ( .IN1(data1[8]), .IN2(n5), .IN3(data0[8]), .IN4(n4), .Q(data_o[8]) );
  AO22X1 U6 ( .IN1(data1[7]), .IN2(n5), .IN3(data0[7]), .IN4(n4), .Q(data_o[7]) );
  AO22X1 U7 ( .IN1(data1[6]), .IN2(n5), .IN3(data0[6]), .IN4(n4), .Q(data_o[6]) );
  AO22X1 U8 ( .IN1(data1[5]), .IN2(n5), .IN3(data0[5]), .IN4(n4), .Q(data_o[5]) );
  AO22X1 U9 ( .IN1(data1[4]), .IN2(n5), .IN3(data0[4]), .IN4(n4), .Q(data_o[4]) );
  AO22X1 U10 ( .IN1(data1[3]), .IN2(n5), .IN3(data0[3]), .IN4(n4), .Q(
        data_o[3]) );
  AO22X1 U11 ( .IN1(data1[2]), .IN2(n5), .IN3(data0[2]), .IN4(n4), .Q(
        data_o[2]) );
  AO22X1 U12 ( .IN1(data1[1]), .IN2(n5), .IN3(data0[1]), .IN4(n4), .Q(
        data_o[1]) );
  AO22X1 U13 ( .IN1(data1[15]), .IN2(n5), .IN3(data0[15]), .IN4(n4), .Q(
        data_o[15]) );
  AO22X1 U14 ( .IN1(data1[14]), .IN2(n5), .IN3(data0[14]), .IN4(n4), .Q(
        data_o[14]) );
  AO22X1 U15 ( .IN1(data1[13]), .IN2(n5), .IN3(data0[13]), .IN4(n4), .Q(
        data_o[13]) );
  AO22X1 U16 ( .IN1(data1[12]), .IN2(n5), .IN3(data0[12]), .IN4(n4), .Q(
        data_o[12]) );
  AO22X1 U17 ( .IN1(data1[11]), .IN2(n5), .IN3(data0[11]), .IN4(n4), .Q(
        data_o[11]) );
  AO22X1 U18 ( .IN1(data1[10]), .IN2(n5), .IN3(data0[10]), .IN4(n4), .Q(
        data_o[10]) );
  AO22X1 U19 ( .IN1(data1[0]), .IN2(n5), .IN3(data0[0]), .IN4(n4), .Q(
        data_o[0]) );
  INVX0 U2 ( .INP(select1), .ZN(n1) );
  AND2X1 U3 ( .IN1(select0), .IN2(n1), .Q(n4) );
  NOR2X0 U20 ( .IN1(n1), .IN2(select0), .QN(n5) );
endmodule


module mux3_1_5 ( data0, data1, data2, select0, select1, select2, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  output [15:0] data_o;
  input select0, select1, select2;
  wire   n1, n2, n6, n7, n8;

  AO222X1 U4 ( .IN1(data1[9]), .IN2(n8), .IN3(data0[9]), .IN4(n7), .IN5(
        data2[9]), .IN6(n6), .Q(data_o[9]) );
  AO222X1 U5 ( .IN1(data1[8]), .IN2(n8), .IN3(data0[8]), .IN4(n7), .IN5(
        data2[8]), .IN6(n6), .Q(data_o[8]) );
  AO222X1 U6 ( .IN1(data1[7]), .IN2(n8), .IN3(data0[7]), .IN4(n7), .IN5(
        data2[7]), .IN6(n6), .Q(data_o[7]) );
  AO222X1 U7 ( .IN1(data1[6]), .IN2(n8), .IN3(data0[6]), .IN4(n7), .IN5(
        data2[6]), .IN6(n6), .Q(data_o[6]) );
  AO222X1 U8 ( .IN1(data1[5]), .IN2(n8), .IN3(data0[5]), .IN4(n7), .IN5(
        data2[5]), .IN6(n6), .Q(data_o[5]) );
  AO222X1 U9 ( .IN1(data1[4]), .IN2(n8), .IN3(data0[4]), .IN4(n7), .IN5(
        data2[4]), .IN6(n6), .Q(data_o[4]) );
  AO222X1 U10 ( .IN1(data1[3]), .IN2(n8), .IN3(data0[3]), .IN4(n7), .IN5(
        data2[3]), .IN6(n6), .Q(data_o[3]) );
  AO222X1 U11 ( .IN1(data1[2]), .IN2(n8), .IN3(data0[2]), .IN4(n7), .IN5(
        data2[2]), .IN6(n6), .Q(data_o[2]) );
  AO222X1 U12 ( .IN1(data1[1]), .IN2(n8), .IN3(data0[1]), .IN4(n7), .IN5(
        data2[1]), .IN6(n6), .Q(data_o[1]) );
  AO222X1 U13 ( .IN1(data1[15]), .IN2(n8), .IN3(data0[15]), .IN4(n7), .IN5(
        data2[15]), .IN6(n6), .Q(data_o[15]) );
  AO222X1 U14 ( .IN1(data1[14]), .IN2(n8), .IN3(data0[14]), .IN4(n7), .IN5(
        data2[14]), .IN6(n6), .Q(data_o[14]) );
  AO222X1 U15 ( .IN1(data1[13]), .IN2(n8), .IN3(data0[13]), .IN4(n7), .IN5(
        data2[13]), .IN6(n6), .Q(data_o[13]) );
  AO222X1 U16 ( .IN1(data1[12]), .IN2(n8), .IN3(data0[12]), .IN4(n7), .IN5(
        data2[12]), .IN6(n6), .Q(data_o[12]) );
  AO222X1 U17 ( .IN1(data1[11]), .IN2(n8), .IN3(data0[11]), .IN4(n7), .IN5(
        data2[11]), .IN6(n6), .Q(data_o[11]) );
  AO222X1 U18 ( .IN1(data1[10]), .IN2(n8), .IN3(data0[10]), .IN4(n7), .IN5(
        data2[10]), .IN6(n6), .Q(data_o[10]) );
  AO222X1 U19 ( .IN1(data1[0]), .IN2(n8), .IN3(data0[0]), .IN4(n7), .IN5(
        data2[0]), .IN6(n6), .Q(data_o[0]) );
  INVX0 U2 ( .INP(select0), .ZN(n2) );
  INVX0 U3 ( .INP(select1), .ZN(n1) );
  AND3X1 U20 ( .IN1(n2), .IN2(n1), .IN3(select2), .Q(n6) );
  NOR3X0 U21 ( .IN1(select1), .IN2(select2), .IN3(n2), .QN(n7) );
  NOR3X0 U22 ( .IN1(select0), .IN2(select2), .IN3(n1), .QN(n8) );
endmodule


module mux3_1_4 ( data0, data1, data2, select0, select1, select2, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  output [15:0] data_o;
  input select0, select1, select2;
  wire   n1, n2, n6, n7, n8;

  AO222X1 U4 ( .IN1(data1[9]), .IN2(n8), .IN3(data0[9]), .IN4(n7), .IN5(
        data2[9]), .IN6(n6), .Q(data_o[9]) );
  AO222X1 U5 ( .IN1(data1[8]), .IN2(n8), .IN3(data0[8]), .IN4(n7), .IN5(
        data2[8]), .IN6(n6), .Q(data_o[8]) );
  AO222X1 U6 ( .IN1(data1[7]), .IN2(n8), .IN3(data0[7]), .IN4(n7), .IN5(
        data2[7]), .IN6(n6), .Q(data_o[7]) );
  AO222X1 U7 ( .IN1(data1[6]), .IN2(n8), .IN3(data0[6]), .IN4(n7), .IN5(
        data2[6]), .IN6(n6), .Q(data_o[6]) );
  AO222X1 U8 ( .IN1(data1[5]), .IN2(n8), .IN3(data0[5]), .IN4(n7), .IN5(
        data2[5]), .IN6(n6), .Q(data_o[5]) );
  AO222X1 U9 ( .IN1(data1[4]), .IN2(n8), .IN3(data0[4]), .IN4(n7), .IN5(
        data2[4]), .IN6(n6), .Q(data_o[4]) );
  AO222X1 U10 ( .IN1(data1[3]), .IN2(n8), .IN3(data0[3]), .IN4(n7), .IN5(
        data2[3]), .IN6(n6), .Q(data_o[3]) );
  AO222X1 U11 ( .IN1(data1[2]), .IN2(n8), .IN3(data0[2]), .IN4(n7), .IN5(
        data2[2]), .IN6(n6), .Q(data_o[2]) );
  AO222X1 U12 ( .IN1(data1[1]), .IN2(n8), .IN3(data0[1]), .IN4(n7), .IN5(
        data2[1]), .IN6(n6), .Q(data_o[1]) );
  AO222X1 U13 ( .IN1(data1[15]), .IN2(n8), .IN3(data0[15]), .IN4(n7), .IN5(
        data2[15]), .IN6(n6), .Q(data_o[15]) );
  AO222X1 U14 ( .IN1(data1[14]), .IN2(n8), .IN3(data0[14]), .IN4(n7), .IN5(
        data2[14]), .IN6(n6), .Q(data_o[14]) );
  AO222X1 U15 ( .IN1(data1[13]), .IN2(n8), .IN3(data0[13]), .IN4(n7), .IN5(
        data2[13]), .IN6(n6), .Q(data_o[13]) );
  AO222X1 U16 ( .IN1(data1[12]), .IN2(n8), .IN3(data0[12]), .IN4(n7), .IN5(
        data2[12]), .IN6(n6), .Q(data_o[12]) );
  AO222X1 U17 ( .IN1(data1[11]), .IN2(n8), .IN3(data0[11]), .IN4(n7), .IN5(
        data2[11]), .IN6(n6), .Q(data_o[11]) );
  AO222X1 U18 ( .IN1(data1[10]), .IN2(n8), .IN3(data0[10]), .IN4(n7), .IN5(
        data2[10]), .IN6(n6), .Q(data_o[10]) );
  AO222X1 U19 ( .IN1(data1[0]), .IN2(n8), .IN3(data0[0]), .IN4(n7), .IN5(
        data2[0]), .IN6(n6), .Q(data_o[0]) );
  INVX0 U2 ( .INP(select0), .ZN(n2) );
  INVX0 U3 ( .INP(select1), .ZN(n1) );
  AND3X1 U20 ( .IN1(n2), .IN2(n1), .IN3(select2), .Q(n6) );
  NOR3X0 U21 ( .IN1(select1), .IN2(select2), .IN3(n2), .QN(n7) );
  NOR3X0 U22 ( .IN1(select0), .IN2(select2), .IN3(n1), .QN(n8) );
endmodule



    module node4_NODE_X0_NODE_Y2I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__I_node_2_node_interface__ ( 
        \clk.clk , \reset.reset , \local_node.clk , 
        \local_node.buffer_full_in , \local_node.buffer_full_out , 
        \local_node.receiving_data , \local_node.sending_data , 
        \local_node.data_in , \local_node.data_out , \node_0.clk , 
        \node_0.buffer_full_in , \node_0.buffer_full_out , 
        \node_0.receiving_data , \node_0.sending_data , \node_0.data_in , 
        \node_0.data_out , \node_1.clk , \node_1.buffer_full_in , 
        \node_1.buffer_full_out , \node_1.receiving_data , 
        \node_1.sending_data , \node_1.data_in , \node_1.data_out , 
        \node_2.clk , \node_2.buffer_full_in , \node_2.buffer_full_out , 
        \node_2.receiving_data , \node_2.sending_data , \node_2.data_in , 
        \node_2.data_out  );
  input [15:0] \local_node.data_in ;
  output [15:0] \local_node.data_out ;
  input [15:0] \node_0.data_in ;
  output [15:0] \node_0.data_out ;
  input [15:0] \node_1.data_in ;
  output [15:0] \node_1.data_out ;
  input [15:0] \node_2.data_in ;
  output [15:0] \node_2.data_out ;
  input \clk.clk , \reset.reset , \local_node.buffer_full_in ,
         \local_node.receiving_data , \node_0.buffer_full_in ,
         \node_0.receiving_data , \node_1.buffer_full_in ,
         \node_1.receiving_data , \node_2.buffer_full_in ,
         \node_2.receiving_data ;
  output \local_node.buffer_full_out , \local_node.sending_data ,
         \node_0.buffer_full_out , \node_0.sending_data ,
         \node_1.buffer_full_out , \node_1.sending_data ,
         \node_2.buffer_full_out , \node_2.sending_data ;
  inout \local_node.clk ,  \node_0.clk ,  \node_1.clk ,  \node_2.clk ;
  wire   \buffer_out[3][15] , \buffer_out[3][14] , \buffer_out[3][13] ,
         \buffer_out[3][12] , \buffer_out[3][11] , \buffer_out[3][10] ,
         \buffer_out[3][9] , \buffer_out[3][8] , \buffer_out[3][7] ,
         \buffer_out[3][6] , \buffer_out[3][5] , \buffer_out[3][4] ,
         \buffer_out[3][3] , \buffer_out[3][2] , \buffer_out[3][1] ,
         \buffer_out[3][0] , \buffer_out[2][15] , \buffer_out[2][14] ,
         \buffer_out[2][13] , \buffer_out[2][12] , \buffer_out[2][11] ,
         \buffer_out[2][10] , \buffer_out[2][9] , \buffer_out[2][8] ,
         \buffer_out[2][7] , \buffer_out[2][6] , \buffer_out[2][5] ,
         \buffer_out[2][4] , \buffer_out[2][3] , \buffer_out[2][2] ,
         \buffer_out[2][1] , \buffer_out[2][0] , \buffer_out[1][15] ,
         \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] ,
         \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] ,
         \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] ,
         \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] ,
         \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] ,
         \buffer_out[0][15] , \buffer_out[0][14] , \buffer_out[0][13] ,
         \buffer_out[0][12] , \buffer_out[0][11] , \buffer_out[0][10] ,
         \buffer_out[0][9] , \buffer_out[0][8] , \buffer_out[0][7] ,
         \buffer_out[0][6] , \buffer_out[0][5] , \buffer_out[0][4] ,
         \buffer_out[0][3] , \buffer_out[0][2] , \buffer_out[0][1] ,
         \buffer_out[0][0] , \next_buffer_out[3][15] ,
         \next_buffer_out[3][14] , \next_buffer_out[3][13] ,
         \next_buffer_out[3][12] , \next_buffer_out[3][11] ,
         \next_buffer_out[3][10] , \next_buffer_out[3][9] ,
         \next_buffer_out[3][8] , \next_buffer_out[3][7] ,
         \next_buffer_out[3][6] , \next_buffer_out[3][5] ,
         \next_buffer_out[3][4] , \next_buffer_out[3][3] ,
         \next_buffer_out[3][2] , \next_buffer_out[3][1] ,
         \next_buffer_out[3][0] , \next_buffer_out[2][15] ,
         \next_buffer_out[2][14] , \next_buffer_out[2][13] ,
         \next_buffer_out[2][12] , \next_buffer_out[2][11] ,
         \next_buffer_out[2][10] , \next_buffer_out[2][9] ,
         \next_buffer_out[2][8] , \next_buffer_out[2][7] ,
         \next_buffer_out[2][6] , \next_buffer_out[2][5] ,
         \next_buffer_out[2][4] , \next_buffer_out[2][3] ,
         \next_buffer_out[2][2] , \next_buffer_out[2][1] ,
         \next_buffer_out[2][0] , \next_buffer_out[1][15] ,
         \next_buffer_out[1][14] , \next_buffer_out[1][13] ,
         \next_buffer_out[1][12] , \next_buffer_out[1][11] ,
         \next_buffer_out[1][10] , \next_buffer_out[1][9] ,
         \next_buffer_out[1][8] , \next_buffer_out[1][7] ,
         \next_buffer_out[1][6] , \next_buffer_out[1][5] ,
         \next_buffer_out[1][4] , \next_buffer_out[1][3] ,
         \next_buffer_out[1][2] , \next_buffer_out[1][1] ,
         \next_buffer_out[1][0] , \next_buffer_out[0][15] ,
         \next_buffer_out[0][14] , \next_buffer_out[0][13] ,
         \next_buffer_out[0][12] , \next_buffer_out[0][11] ,
         \next_buffer_out[0][10] , \next_buffer_out[0][9] ,
         \next_buffer_out[0][8] , \next_buffer_out[0][7] ,
         \next_buffer_out[0][6] , \next_buffer_out[0][5] ,
         \next_buffer_out[0][4] , \next_buffer_out[0][3] ,
         \next_buffer_out[0][2] , \next_buffer_out[0][1] ,
         \next_buffer_out[0][0] ;
  wire   [3:0] buffer_full_in;
  wire   [3:0] receiving_data;
  wire   [3:0] pop_v;
  wire   [3:0] data_valid;
  wire   [3:0] next_data_valid;
  wire   [1:0] grant_0;
  wire   [1:0] grant_1;
  wire   [2:0] grant_2;
  wire   [2:0] grant_3;
  tri   \local_node.buffer_full_in ;
  tri   \local_node.buffer_full_out ;
  tri   \local_node.receiving_data ;
  tri   \local_node.sending_data ;
  tri   [15:0] \local_node.data_in ;
  tri   [15:0] \local_node.data_out ;

  converter_out_I_n_node_interface_dut_ c3 ( .\n.buffer_full_in (
        \local_node.buffer_full_in ), .\n.receiving_data (
        \local_node.receiving_data ), .\n.data_in (\local_node.data_in ), 
        .\n.buffer_full_out (\local_node.buffer_full_out ), .\n.sending_data (
        \local_node.sending_data ), .\n.data_out (\local_node.data_out ), 
        .buffer_full_in(1'b0), .receiving_data(1'b0), .data_in({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  fifo_kev_31 \genblk1[0].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[0]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[0]), .data_out({\buffer_out[0][15] , 
        \buffer_out[0][14] , \buffer_out[0][13] , \buffer_out[0][12] , 
        \buffer_out[0][11] , \buffer_out[0][10] , \buffer_out[0][9] , 
        \buffer_out[0][8] , \buffer_out[0][7] , \buffer_out[0][6] , 
        \buffer_out[0][5] , \buffer_out[0][4] , \buffer_out[0][3] , 
        \buffer_out[0][2] , \buffer_out[0][1] , \buffer_out[0][0] }), 
        .next_data_out({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] , 
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .next_data_valid(
        next_data_valid[0]) );
  address_counter_31 \genblk1[0].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] }), 
        .buffer_data_valid(next_data_valid[0]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .buffer_pop(
        pop_v[0]), .receiving_data(1'b0) );
  fifo_kev_30 \genblk1[1].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[1]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[1]), .data_out({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), 
        .next_data_out({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] , 
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .next_data_valid(
        next_data_valid[1]) );
  address_counter_30 \genblk1[1].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] }), 
        .buffer_data_valid(next_data_valid[1]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .buffer_pop(
        pop_v[1]), .receiving_data(1'b0) );
  fifo_kev_29 \genblk1[2].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[2]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[2]), .data_out({\buffer_out[2][15] , 
        \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] , 
        \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] , 
        \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] , 
        \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] , 
        \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] }), 
        .next_data_out({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] , 
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .next_data_valid(
        next_data_valid[2]) );
  address_counter_29 \genblk1[2].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] }), 
        .buffer_data_valid(next_data_valid[2]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .buffer_pop(
        pop_v[2]), .receiving_data(1'b0) );
  fifo_kev_28 \genblk1[3].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[3]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[3]), .data_out({\buffer_out[3][15] , 
        \buffer_out[3][14] , \buffer_out[3][13] , \buffer_out[3][12] , 
        \buffer_out[3][11] , \buffer_out[3][10] , \buffer_out[3][9] , 
        \buffer_out[3][8] , \buffer_out[3][7] , \buffer_out[3][6] , 
        \buffer_out[3][5] , \buffer_out[3][4] , \buffer_out[3][3] , 
        \buffer_out[3][2] , \buffer_out[3][1] , \buffer_out[3][0] }), 
        .next_data_out({\next_buffer_out[3][15] , \next_buffer_out[3][14] , 
        \next_buffer_out[3][13] , \next_buffer_out[3][12] , 
        \next_buffer_out[3][11] , \next_buffer_out[3][10] , 
        \next_buffer_out[3][9] , \next_buffer_out[3][8] , 
        \next_buffer_out[3][7] , \next_buffer_out[3][6] , 
        \next_buffer_out[3][5] , \next_buffer_out[3][4] , 
        \next_buffer_out[3][3] , \next_buffer_out[3][2] , 
        \next_buffer_out[3][1] , \next_buffer_out[3][0] }), .next_data_valid(
        next_data_valid[3]) );
  address_counter_28 \genblk1[3].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[3][15] , \next_buffer_out[3][14] , 
        \next_buffer_out[3][13] , \next_buffer_out[3][12] , 
        \next_buffer_out[3][11] , \next_buffer_out[3][10] , 
        \next_buffer_out[3][9] , \next_buffer_out[3][8] }), 
        .buffer_data_valid(next_data_valid[3]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[3][7] , \next_buffer_out[3][6] , 
        \next_buffer_out[3][5] , \next_buffer_out[3][4] , 
        \next_buffer_out[3][3] , \next_buffer_out[3][2] , 
        \next_buffer_out[3][1] , \next_buffer_out[3][0] }), .buffer_pop(
        pop_v[3]), .receiving_data(1'b0) );
  converter_in_I_n_node_interface_dut__11 \genblk2.c0  ( .\n.buffer_full_in (
        \node_0.buffer_full_in ), .\n.receiving_data (\node_0.receiving_data ), 
        .\n.data_in (\node_0.data_in ), .\n.buffer_full_out (
        \node_0.buffer_full_out ), .\n.sending_data (\node_0.sending_data ), 
        .\n.data_out (\node_0.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_out_I_n_node_interface_dut_ \genblk2.c1  ( .\n.buffer_full_in (
        \node_1.buffer_full_in ), .\n.receiving_data (\node_1.receiving_data ), 
        .\n.data_in (\node_1.data_in ), .\n.buffer_full_out (
        \node_1.buffer_full_out ), .\n.sending_data (\node_1.sending_data ), 
        .\n.data_out (\node_1.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_in_I_n_node_interface_dut__10 \genblk2.c2  ( .\n.buffer_full_in (
        \node_2.buffer_full_in ), .\n.receiving_data (\node_2.receiving_data ), 
        .\n.data_in (\node_2.data_in ), .\n.buffer_full_out (
        \node_2.buffer_full_out ), .\n.sending_data (\node_2.sending_data ), 
        .\n.data_out (\node_2.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  controller4_edge_w_0 \genblk2.w  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .packet_addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .local_addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0}), 
        .packet_valid(data_valid), .buffer_full_in({1'b0, 1'b0, 1'b0, 1'b0}), 
        .grant_0(grant_0), .grant_1(grant_1), .grant_2(grant_2), .grant_3(
        grant_3), .pop_v(pop_v) );
  mux2_1_13 \genblk2.mux_n  ( .data0({\buffer_out[1][15] , \buffer_out[1][14] , 
        \buffer_out[1][13] , \buffer_out[1][12] , \buffer_out[1][11] , 
        \buffer_out[1][10] , \buffer_out[1][9] , \buffer_out[1][8] , 
        \buffer_out[1][7] , \buffer_out[1][6] , \buffer_out[1][5] , 
        \buffer_out[1][4] , \buffer_out[1][3] , \buffer_out[1][2] , 
        \buffer_out[1][1] , \buffer_out[1][0] }), .data1({\buffer_out[3][15] , 
        \buffer_out[3][14] , \buffer_out[3][13] , \buffer_out[3][12] , 
        \buffer_out[3][11] , \buffer_out[3][10] , \buffer_out[3][9] , 
        \buffer_out[3][8] , \buffer_out[3][7] , \buffer_out[3][6] , 
        \buffer_out[3][5] , \buffer_out[3][4] , \buffer_out[3][3] , 
        \buffer_out[3][2] , \buffer_out[3][1] , \buffer_out[3][0] }), 
        .select0(grant_0[0]), .select1(grant_0[1]) );
  mux2_1_12 \genblk2.mux_s  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[3][15] , 
        \buffer_out[3][14] , \buffer_out[3][13] , \buffer_out[3][12] , 
        \buffer_out[3][11] , \buffer_out[3][10] , \buffer_out[3][9] , 
        \buffer_out[3][8] , \buffer_out[3][7] , \buffer_out[3][6] , 
        \buffer_out[3][5] , \buffer_out[3][4] , \buffer_out[3][3] , 
        \buffer_out[3][2] , \buffer_out[3][1] , \buffer_out[3][0] }), 
        .select0(grant_1[0]), .select1(grant_1[1]) );
  mux3_1_5 \genblk2.mux_e  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[3][15] , \buffer_out[3][14] , \buffer_out[3][13] , 
        \buffer_out[3][12] , \buffer_out[3][11] , \buffer_out[3][10] , 
        \buffer_out[3][9] , \buffer_out[3][8] , \buffer_out[3][7] , 
        \buffer_out[3][6] , \buffer_out[3][5] , \buffer_out[3][4] , 
        \buffer_out[3][3] , \buffer_out[3][2] , \buffer_out[3][1] , 
        \buffer_out[3][0] }), .select0(grant_2[0]), .select1(grant_2[1]), 
        .select2(grant_2[2]) );
  mux3_1_4 \genblk2.mux_l  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[2][15] , \buffer_out[2][14] , \buffer_out[2][13] , 
        \buffer_out[2][12] , \buffer_out[2][11] , \buffer_out[2][10] , 
        \buffer_out[2][9] , \buffer_out[2][8] , \buffer_out[2][7] , 
        \buffer_out[2][6] , \buffer_out[2][5] , \buffer_out[2][4] , 
        \buffer_out[2][3] , \buffer_out[2][2] , \buffer_out[2][1] , 
        \buffer_out[2][0] }), .select0(grant_3[0]), .select1(grant_3[1]), 
        .select2(grant_3[2]) );
endmodule


module fifo_kev_27 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_55 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_27 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_55 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_54 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_27 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_54 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_27_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_27 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_27 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_27 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_27_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_26 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_53 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_26 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_53 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_52 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_26 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_52 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_26_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_26 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_26 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_26 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_26_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_25 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_51 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_25 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_51 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_50 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_25 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_50 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_25_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_25 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_25 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_25 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_25_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_24 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_49 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_24 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_49 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_48 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_24 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_48 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_24_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_24 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_24 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_24 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_24_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module converter_in_I_n_node_interface_dut__9 ( \n.buffer_full_in , 
        \n.receiving_data , \n.data_in , \n.buffer_full_out , \n.sending_data , 
        \n.data_out , buffer_full_out, sending_data, data_out, buffer_full_in, 
        receiving_data, data_in );
  input [15:0] \n.data_in ;
  output [15:0] \n.data_out ;
  output [15:0] data_out;
  input [15:0] data_in;
  input \n.buffer_full_in , \n.receiving_data , buffer_full_in, receiving_data;
  output \n.buffer_full_out , \n.sending_data , buffer_full_out, sending_data;
  wire   \n.buffer_full_in , \n.receiving_data , buffer_full_in,
         receiving_data;
  assign buffer_full_out = \n.buffer_full_in ;
  assign sending_data = \n.receiving_data ;
  assign data_out[15] = \n.data_in  [15];
  assign data_out[14] = \n.data_in  [14];
  assign data_out[13] = \n.data_in  [13];
  assign data_out[12] = \n.data_in  [12];
  assign data_out[11] = \n.data_in  [11];
  assign data_out[10] = \n.data_in  [10];
  assign data_out[9] = \n.data_in  [9];
  assign data_out[8] = \n.data_in  [8];
  assign data_out[7] = \n.data_in  [7];
  assign data_out[6] = \n.data_in  [6];
  assign data_out[5] = \n.data_in  [5];
  assign data_out[4] = \n.data_in  [4];
  assign data_out[3] = \n.data_in  [3];
  assign data_out[2] = \n.data_in  [2];
  assign data_out[1] = \n.data_in  [1];
  assign data_out[0] = \n.data_in  [0];
  assign \n.buffer_full_out  = buffer_full_in;
  assign \n.sending_data  = receiving_data;
  assign \n.data_out  [15] = data_in[15];
  assign \n.data_out  [14] = data_in[14];
  assign \n.data_out  [13] = data_in[13];
  assign \n.data_out  [12] = data_in[12];
  assign \n.data_out  [11] = data_in[11];
  assign \n.data_out  [10] = data_in[10];
  assign \n.data_out  [9] = data_in[9];
  assign \n.data_out  [8] = data_in[8];
  assign \n.data_out  [7] = data_in[7];
  assign \n.data_out  [6] = data_in[6];
  assign \n.data_out  [5] = data_in[5];
  assign \n.data_out  [4] = data_in[4];
  assign \n.data_out  [3] = data_in[3];
  assign \n.data_out  [2] = data_in[2];
  assign \n.data_out  [1] = data_in[1];
  assign \n.data_out  [0] = data_in[0];

endmodule


module flipflop_BITS2_11 ( clk, data_i, data_o );
  input [1:0] data_i;
  output [1:0] data_o;
  input clk;


  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS2_11 ( clk, enable_i, reset, data_i, data_o );
  input [1:0] data_i;
  input [1:0] data_o;
  input clk, enable_i, reset;
  wire   n10, n11, n1, n5, n7, n8, n9;
  wire   [1:0] write_data;

  AOI22X1 U5 ( .IN1(enable_i), .IN2(data_i[1]), .IN3(n10), .IN4(n1), .QN(n9)
         );
  AOI22X1 U6 ( .IN1(data_i[0]), .IN2(enable_i), .IN3(n11), .IN4(n1), .QN(n8)
         );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n9), .QN(write_data[1]) );
  NOR2X0 U4 ( .IN1(reset), .IN2(n8), .QN(write_data[0]) );
  AND2X1 U7 ( .IN1(data_o[1]), .IN2(n7), .Q(n10) );
  AND2X1 U8 ( .IN1(data_o[0]), .IN2(n5), .Q(n11) );
  flipflop_BITS2_11 FF ( .clk(clk), .data_i(write_data), .data_o({n7, n5}) );
endmodule


module flipflop_BITS1_43 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_43 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_43 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter2_11 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [1:0] request;
  output [1:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   tail_en, n1, n2;
  wire   [1:0] req_i;
  wire   [1:0] req_o;

  AND3X1 U10 ( .IN1(request[1]), .IN2(n1), .IN3(n2), .Q(grant[1]) );
  AND3X1 U11 ( .IN1(request[0]), .IN2(n2), .IN3(request[1]), .Q(tail_en) );
  INVX0 U6 ( .INP(request[0]), .ZN(n1) );
  NOR2X0 U7 ( .IN1(buffer_full_i), .IN2(n1), .QN(grant[0]) );
  INVX0 U8 ( .INP(buffer_full_i), .ZN(n2) );
  OA21X1 U9 ( .IN1(request[1]), .IN2(request[0]), .IN3(n2), .Q(grant_v_o) );
  register_BITS2_11 req_record ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i({1'b1, 1'b0}), .data_o({1'b0, 1'b0}) );
  register_BITS1_43 tail ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i(1'b1), .data_o(1'b0) );
endmodule


module flipflop_BITS2_10 ( clk, data_i, data_o );
  input [1:0] data_i;
  output [1:0] data_o;
  input clk;


  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS2_10 ( clk, enable_i, reset, data_i, data_o );
  input [1:0] data_i;
  input [1:0] data_o;
  input clk, enable_i, reset;
  wire   n10, n11, n1, n5, n7, n8, n9;
  wire   [1:0] write_data;

  AOI22X1 U5 ( .IN1(enable_i), .IN2(data_i[1]), .IN3(n10), .IN4(n1), .QN(n9)
         );
  AOI22X1 U6 ( .IN1(data_i[0]), .IN2(enable_i), .IN3(n11), .IN4(n1), .QN(n8)
         );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n9), .QN(write_data[1]) );
  NOR2X0 U4 ( .IN1(reset), .IN2(n8), .QN(write_data[0]) );
  AND2X1 U7 ( .IN1(data_o[1]), .IN2(n7), .Q(n10) );
  AND2X1 U8 ( .IN1(data_o[0]), .IN2(n5), .Q(n11) );
  flipflop_BITS2_10 FF ( .clk(clk), .data_i(write_data), .data_o({n7, n5}) );
endmodule


module flipflop_BITS1_42 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_42 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_42 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter2_10 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [1:0] request;
  output [1:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   tail_en, n1, n2;
  wire   [1:0] req_i;
  wire   [1:0] req_o;

  AND3X1 U10 ( .IN1(request[1]), .IN2(n1), .IN3(n2), .Q(grant[1]) );
  AND3X1 U11 ( .IN1(request[0]), .IN2(n2), .IN3(request[1]), .Q(tail_en) );
  INVX0 U6 ( .INP(request[0]), .ZN(n1) );
  NOR2X0 U7 ( .IN1(buffer_full_i), .IN2(n1), .QN(grant[0]) );
  INVX0 U8 ( .INP(buffer_full_i), .ZN(n2) );
  OA21X1 U9 ( .IN1(request[1]), .IN2(request[0]), .IN3(n2), .Q(grant_v_o) );
  register_BITS2_10 req_record ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i({1'b1, 1'b0}), .data_o({1'b0, 1'b0}) );
  register_BITS1_42 tail ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i(1'b1), .data_o(1'b0) );
endmodule


module flipflop_BITS3_7 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_7 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_7 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS3_6 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_6 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_6 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS1_41 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_41 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_41 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_40 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_40 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_40 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter3_3 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [2:0] request;
  output [2:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[1][2] , \req_i[1][1] , \req_i[1][0] , \req_i[0][2] ,
         \req_i[0][1] , tail_en, N99, N100, N101, N110, N111, N118, N119, N120,
         N121, n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [1:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N99 = request[0];
  assign N100 = request[1];
  assign N101 = request[2];

  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(N111), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(N110), .Q(\req_i[0][1] ) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N121), .D(tail_en), .Q(req_en[0]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N120), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N119), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N118), .Q(grant[0]) );
  AND2X1 U20 ( .IN1(n8), .IN2(N101), .Q(n7) );
  OR3X1 U21 ( .IN1(n3), .IN2(N111), .IN3(n6), .Q(N121) );
  NOR3X0 U22 ( .IN1(N99), .IN2(N100), .IN3(n6), .QN(N120) );
  NOR3X0 U23 ( .IN1(n2), .IN2(N99), .IN3(n6), .QN(N119) );
  NAND3X0 U24 ( .IN1(n2), .IN2(n3), .IN3(n1), .QN(n5) );
  AO22X1 U25 ( .IN1(N100), .IN2(N101), .IN3(N99), .IN4(N101), .Q(N111) );
  INVX0 U10 ( .INP(N101), .ZN(n3) );
  NAND2X1 U11 ( .IN1(n5), .IN2(n4), .QN(n6) );
  INVX0 U12 ( .INP(N99), .ZN(n1) );
  INVX0 U13 ( .INP(N100), .ZN(n2) );
  INVX0 U14 ( .INP(buffer_full_i), .ZN(n4) );
  NAND2X1 U15 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NOR2X0 U16 ( .IN1(n1), .IN2(n6), .QN(N118) );
  NOR2X0 U17 ( .IN1(n1), .IN2(n2), .QN(N110) );
  OA21X1 U18 ( .IN1(N110), .IN2(n7), .IN3(n4), .Q(tail_en) );
  OA21X1 U19 ( .IN1(N101), .IN2(n8), .IN3(n4), .Q(grant_v_o) );
  register_BITS3_7 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][2] , \req_i[0][1] , 1'b0}), .data_o({
        1'b0, 1'b0, 1'b0}) );
  register_BITS3_6 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][2] , \req_i[1][1] , \req_i[1][0] }), 
        .data_o({1'b0, 1'b0, 1'b0}) );
  register_BITS1_41 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b1), .data_o(1'b0) );
  register_BITS1_40 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module flipflop_BITS3_5 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_5 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_5 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS3_4 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_4 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_4 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS1_39 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_39 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_39 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_38 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_38 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_38 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter3_2 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [2:0] request;
  output [2:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[1][2] , \req_i[1][1] , \req_i[1][0] , \req_i[0][2] ,
         \req_i[0][1] , tail_en, N99, N100, N101, N110, N111, N118, N119, N120,
         N121, n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [1:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N99 = request[0];
  assign N100 = request[1];
  assign N101 = request[2];

  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(N111), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(N110), .Q(\req_i[0][1] ) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N121), .D(tail_en), .Q(req_en[0]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N120), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N119), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N118), .Q(grant[0]) );
  AND2X1 U20 ( .IN1(n8), .IN2(N101), .Q(n7) );
  OR3X1 U21 ( .IN1(n3), .IN2(N111), .IN3(n6), .Q(N121) );
  NOR3X0 U22 ( .IN1(N99), .IN2(N100), .IN3(n6), .QN(N120) );
  NOR3X0 U23 ( .IN1(n2), .IN2(N99), .IN3(n6), .QN(N119) );
  NAND3X0 U24 ( .IN1(n2), .IN2(n3), .IN3(n1), .QN(n5) );
  AO22X1 U25 ( .IN1(N100), .IN2(N101), .IN3(N99), .IN4(N101), .Q(N111) );
  INVX0 U10 ( .INP(N101), .ZN(n3) );
  NAND2X1 U11 ( .IN1(n5), .IN2(n4), .QN(n6) );
  INVX0 U12 ( .INP(N99), .ZN(n1) );
  INVX0 U13 ( .INP(N100), .ZN(n2) );
  INVX0 U14 ( .INP(buffer_full_i), .ZN(n4) );
  NAND2X1 U15 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NOR2X0 U16 ( .IN1(n1), .IN2(n6), .QN(N118) );
  NOR2X0 U17 ( .IN1(n1), .IN2(n2), .QN(N110) );
  OA21X1 U18 ( .IN1(N110), .IN2(n7), .IN3(n4), .Q(tail_en) );
  OA21X1 U19 ( .IN1(N101), .IN2(n8), .IN3(n4), .Q(grant_v_o) );
  register_BITS3_5 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][2] , \req_i[0][1] , 1'b0}), .data_o({
        1'b0, 1'b0, 1'b0}) );
  register_BITS3_4 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][2] , \req_i[1][1] , \req_i[1][0] }), 
        .data_o({1'b0, 1'b0, 1'b0}) );
  register_BITS1_39 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b1), .data_o(1'b0) );
  register_BITS1_38 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module dccl_27 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_26 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_25 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_24 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module controller4_edge_e_1 ( clk, rst, .packet_addr({\packet_addr[3][7] , 
        \packet_addr[3][6] , \packet_addr[3][5] , \packet_addr[3][4] , 
        \packet_addr[3][3] , \packet_addr[3][2] , \packet_addr[3][1] , 
        \packet_addr[3][0] , \packet_addr[2][7] , \packet_addr[2][6] , 
        \packet_addr[2][5] , \packet_addr[2][4] , \packet_addr[2][3] , 
        \packet_addr[2][2] , \packet_addr[2][1] , \packet_addr[2][0] , 
        \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] , 
        \packet_addr[1][4] , \packet_addr[1][3] , \packet_addr[1][2] , 
        \packet_addr[1][1] , \packet_addr[1][0] , \packet_addr[0][7] , 
        \packet_addr[0][6] , \packet_addr[0][5] , \packet_addr[0][4] , 
        \packet_addr[0][3] , \packet_addr[0][2] , \packet_addr[0][1] , 
        \packet_addr[0][0] }), local_addr, packet_valid, buffer_full_in, 
        grant_0, grant_1, grant_2, grant_3, grant_v, pop_v );
  input [7:0] local_addr;
  input [3:0] packet_valid;
  input [3:0] buffer_full_in;
  output [1:0] grant_0;
  output [1:0] grant_1;
  output [2:0] grant_2;
  output [2:0] grant_3;
  output [3:0] grant_v;
  output [3:0] pop_v;
  input clk, rst, \packet_addr[3][7] , \packet_addr[3][6] ,
         \packet_addr[3][5] , \packet_addr[3][4] , \packet_addr[3][3] ,
         \packet_addr[3][2] , \packet_addr[3][1] , \packet_addr[3][0] ,
         \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] ,
         \packet_addr[2][4] , \packet_addr[2][3] , \packet_addr[2][2] ,
         \packet_addr[2][1] , \packet_addr[2][0] , \packet_addr[1][7] ,
         \packet_addr[1][6] , \packet_addr[1][5] , \packet_addr[1][4] ,
         \packet_addr[1][3] , \packet_addr[1][2] , \packet_addr[1][1] ,
         \packet_addr[1][0] , \packet_addr[0][7] , \packet_addr[0][6] ,
         \packet_addr[0][5] , \packet_addr[0][4] , \packet_addr[0][3] ,
         \packet_addr[0][2] , \packet_addr[0][1] , \packet_addr[0][0] ;
  wire   \grant_3[2] , \request[3][2] , \request[3][1] , \request[3][0] ,
         \request[2][2] , \request[2][1] , \request[2][0] , \request[1][1] ,
         \request[1][0] , \request[0][1] , \request[0][0] ;
  assign pop_v[2] = \grant_3[2] ;
  assign grant_3[2] = \grant_3[2] ;

  OR3X1 U1 ( .IN1(grant_2[2]), .IN2(grant_1[1]), .IN3(grant_0[1]), .Q(pop_v[3]) );
  OR3X1 U2 ( .IN1(grant_3[1]), .IN2(grant_2[1]), .IN3(grant_0[0]), .Q(pop_v[1]) );
  OR3X1 U3 ( .IN1(grant_3[0]), .IN2(grant_2[0]), .IN3(grant_1[0]), .Q(pop_v[0]) );
  arbiter2_11 arbiter_n ( .clk(clk), .rst(rst), .request({\request[0][1] , 
        \request[0][0] }), .buffer_full_i(buffer_full_in[0]), .grant(grant_0), 
        .grant_v_o(grant_v[0]) );
  arbiter2_10 arbiter_s ( .clk(clk), .rst(rst), .request({\request[1][1] , 
        \request[1][0] }), .buffer_full_i(buffer_full_in[1]), .grant(grant_1), 
        .grant_v_o(grant_v[1]) );
  arbiter3_3 arbiter_w ( .clk(clk), .rst(rst), .request({\request[2][2] , 
        \request[2][1] , \request[2][0] }), .buffer_full_i(buffer_full_in[2]), 
        .grant(grant_2), .grant_v_o(grant_v[2]) );
  arbiter3_2 arbiter_l ( .clk(clk), .rst(rst), .request({\request[3][2] , 
        \request[3][1] , \request[3][0] }), .buffer_full_i(buffer_full_in[3]), 
        .grant({\grant_3[2] , grant_3[1:0]}), .grant_v_o(grant_v[3]) );
  dccl_27 dccl_n ( .packet_addr_y_i({\packet_addr[0][3] , \packet_addr[0][2] , 
        \packet_addr[0][1] , \packet_addr[0][0] }), .packet_addr_x_i({
        \packet_addr[0][7] , \packet_addr[0][6] , \packet_addr[0][5] , 
        \packet_addr[0][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[0]), 
        .south_req(\request[1][0] ), .west_req(\request[2][0] ), .local_req(
        \request[3][0] ) );
  dccl_26 dccl_s ( .packet_addr_y_i({\packet_addr[1][3] , \packet_addr[1][2] , 
        \packet_addr[1][1] , \packet_addr[1][0] }), .packet_addr_x_i({
        \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] , 
        \packet_addr[1][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[1]), 
        .north_req(\request[0][0] ), .west_req(\request[2][1] ), .local_req(
        \request[3][1] ) );
  dccl_25 dccl_w ( .packet_addr_y_i({\packet_addr[2][3] , \packet_addr[2][2] , 
        \packet_addr[2][1] , \packet_addr[2][0] }), .packet_addr_x_i({
        \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] , 
        \packet_addr[2][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[2]), 
        .local_req(\request[3][2] ) );
  dccl_24 dccl_l ( .packet_addr_y_i({\packet_addr[3][3] , \packet_addr[3][2] , 
        \packet_addr[3][1] , \packet_addr[3][0] }), .packet_addr_x_i({
        \packet_addr[3][7] , \packet_addr[3][6] , \packet_addr[3][5] , 
        \packet_addr[3][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[3]), 
        .north_req(\request[0][1] ), .south_req(\request[1][1] ), .west_req(
        \request[2][2] ) );
endmodule


module mux2_1_11 ( data0, data1, select0, select1, data_o );
  input [15:0] data0;
  input [15:0] data1;
  output [15:0] data_o;
  input select0, select1;
  wire   n1, n4, n5;

  AO22X1 U4 ( .IN1(data1[9]), .IN2(n5), .IN3(data0[9]), .IN4(n4), .Q(data_o[9]) );
  AO22X1 U5 ( .IN1(data1[8]), .IN2(n5), .IN3(data0[8]), .IN4(n4), .Q(data_o[8]) );
  AO22X1 U6 ( .IN1(data1[7]), .IN2(n5), .IN3(data0[7]), .IN4(n4), .Q(data_o[7]) );
  AO22X1 U7 ( .IN1(data1[6]), .IN2(n5), .IN3(data0[6]), .IN4(n4), .Q(data_o[6]) );
  AO22X1 U8 ( .IN1(data1[5]), .IN2(n5), .IN3(data0[5]), .IN4(n4), .Q(data_o[5]) );
  AO22X1 U9 ( .IN1(data1[4]), .IN2(n5), .IN3(data0[4]), .IN4(n4), .Q(data_o[4]) );
  AO22X1 U10 ( .IN1(data1[3]), .IN2(n5), .IN3(data0[3]), .IN4(n4), .Q(
        data_o[3]) );
  AO22X1 U11 ( .IN1(data1[2]), .IN2(n5), .IN3(data0[2]), .IN4(n4), .Q(
        data_o[2]) );
  AO22X1 U12 ( .IN1(data1[1]), .IN2(n5), .IN3(data0[1]), .IN4(n4), .Q(
        data_o[1]) );
  AO22X1 U13 ( .IN1(data1[15]), .IN2(n5), .IN3(data0[15]), .IN4(n4), .Q(
        data_o[15]) );
  AO22X1 U14 ( .IN1(data1[14]), .IN2(n5), .IN3(data0[14]), .IN4(n4), .Q(
        data_o[14]) );
  AO22X1 U15 ( .IN1(data1[13]), .IN2(n5), .IN3(data0[13]), .IN4(n4), .Q(
        data_o[13]) );
  AO22X1 U16 ( .IN1(data1[12]), .IN2(n5), .IN3(data0[12]), .IN4(n4), .Q(
        data_o[12]) );
  AO22X1 U17 ( .IN1(data1[11]), .IN2(n5), .IN3(data0[11]), .IN4(n4), .Q(
        data_o[11]) );
  AO22X1 U18 ( .IN1(data1[10]), .IN2(n5), .IN3(data0[10]), .IN4(n4), .Q(
        data_o[10]) );
  AO22X1 U19 ( .IN1(data1[0]), .IN2(n5), .IN3(data0[0]), .IN4(n4), .Q(
        data_o[0]) );
  INVX0 U2 ( .INP(select1), .ZN(n1) );
  AND2X1 U3 ( .IN1(select0), .IN2(n1), .Q(n4) );
  NOR2X0 U20 ( .IN1(n1), .IN2(select0), .QN(n5) );
endmodule


module mux2_1_10 ( data0, data1, select0, select1, data_o );
  input [15:0] data0;
  input [15:0] data1;
  output [15:0] data_o;
  input select0, select1;
  wire   n1, n4, n5;

  AO22X1 U4 ( .IN1(data1[9]), .IN2(n5), .IN3(data0[9]), .IN4(n4), .Q(data_o[9]) );
  AO22X1 U5 ( .IN1(data1[8]), .IN2(n5), .IN3(data0[8]), .IN4(n4), .Q(data_o[8]) );
  AO22X1 U6 ( .IN1(data1[7]), .IN2(n5), .IN3(data0[7]), .IN4(n4), .Q(data_o[7]) );
  AO22X1 U7 ( .IN1(data1[6]), .IN2(n5), .IN3(data0[6]), .IN4(n4), .Q(data_o[6]) );
  AO22X1 U8 ( .IN1(data1[5]), .IN2(n5), .IN3(data0[5]), .IN4(n4), .Q(data_o[5]) );
  AO22X1 U9 ( .IN1(data1[4]), .IN2(n5), .IN3(data0[4]), .IN4(n4), .Q(data_o[4]) );
  AO22X1 U10 ( .IN1(data1[3]), .IN2(n5), .IN3(data0[3]), .IN4(n4), .Q(
        data_o[3]) );
  AO22X1 U11 ( .IN1(data1[2]), .IN2(n5), .IN3(data0[2]), .IN4(n4), .Q(
        data_o[2]) );
  AO22X1 U12 ( .IN1(data1[1]), .IN2(n5), .IN3(data0[1]), .IN4(n4), .Q(
        data_o[1]) );
  AO22X1 U13 ( .IN1(data1[15]), .IN2(n5), .IN3(data0[15]), .IN4(n4), .Q(
        data_o[15]) );
  AO22X1 U14 ( .IN1(data1[14]), .IN2(n5), .IN3(data0[14]), .IN4(n4), .Q(
        data_o[14]) );
  AO22X1 U15 ( .IN1(data1[13]), .IN2(n5), .IN3(data0[13]), .IN4(n4), .Q(
        data_o[13]) );
  AO22X1 U16 ( .IN1(data1[12]), .IN2(n5), .IN3(data0[12]), .IN4(n4), .Q(
        data_o[12]) );
  AO22X1 U17 ( .IN1(data1[11]), .IN2(n5), .IN3(data0[11]), .IN4(n4), .Q(
        data_o[11]) );
  AO22X1 U18 ( .IN1(data1[10]), .IN2(n5), .IN3(data0[10]), .IN4(n4), .Q(
        data_o[10]) );
  AO22X1 U19 ( .IN1(data1[0]), .IN2(n5), .IN3(data0[0]), .IN4(n4), .Q(
        data_o[0]) );
  INVX0 U2 ( .INP(select1), .ZN(n1) );
  AND2X1 U3 ( .IN1(select0), .IN2(n1), .Q(n4) );
  NOR2X0 U20 ( .IN1(n1), .IN2(select0), .QN(n5) );
endmodule


module mux3_1_3 ( data0, data1, data2, select0, select1, select2, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  output [15:0] data_o;
  input select0, select1, select2;
  wire   n1, n2, n6, n7, n8;

  AO222X1 U4 ( .IN1(data1[9]), .IN2(n8), .IN3(data0[9]), .IN4(n7), .IN5(
        data2[9]), .IN6(n6), .Q(data_o[9]) );
  AO222X1 U5 ( .IN1(data1[8]), .IN2(n8), .IN3(data0[8]), .IN4(n7), .IN5(
        data2[8]), .IN6(n6), .Q(data_o[8]) );
  AO222X1 U6 ( .IN1(data1[7]), .IN2(n8), .IN3(data0[7]), .IN4(n7), .IN5(
        data2[7]), .IN6(n6), .Q(data_o[7]) );
  AO222X1 U7 ( .IN1(data1[6]), .IN2(n8), .IN3(data0[6]), .IN4(n7), .IN5(
        data2[6]), .IN6(n6), .Q(data_o[6]) );
  AO222X1 U8 ( .IN1(data1[5]), .IN2(n8), .IN3(data0[5]), .IN4(n7), .IN5(
        data2[5]), .IN6(n6), .Q(data_o[5]) );
  AO222X1 U9 ( .IN1(data1[4]), .IN2(n8), .IN3(data0[4]), .IN4(n7), .IN5(
        data2[4]), .IN6(n6), .Q(data_o[4]) );
  AO222X1 U10 ( .IN1(data1[3]), .IN2(n8), .IN3(data0[3]), .IN4(n7), .IN5(
        data2[3]), .IN6(n6), .Q(data_o[3]) );
  AO222X1 U11 ( .IN1(data1[2]), .IN2(n8), .IN3(data0[2]), .IN4(n7), .IN5(
        data2[2]), .IN6(n6), .Q(data_o[2]) );
  AO222X1 U12 ( .IN1(data1[1]), .IN2(n8), .IN3(data0[1]), .IN4(n7), .IN5(
        data2[1]), .IN6(n6), .Q(data_o[1]) );
  AO222X1 U13 ( .IN1(data1[15]), .IN2(n8), .IN3(data0[15]), .IN4(n7), .IN5(
        data2[15]), .IN6(n6), .Q(data_o[15]) );
  AO222X1 U14 ( .IN1(data1[14]), .IN2(n8), .IN3(data0[14]), .IN4(n7), .IN5(
        data2[14]), .IN6(n6), .Q(data_o[14]) );
  AO222X1 U15 ( .IN1(data1[13]), .IN2(n8), .IN3(data0[13]), .IN4(n7), .IN5(
        data2[13]), .IN6(n6), .Q(data_o[13]) );
  AO222X1 U16 ( .IN1(data1[12]), .IN2(n8), .IN3(data0[12]), .IN4(n7), .IN5(
        data2[12]), .IN6(n6), .Q(data_o[12]) );
  AO222X1 U17 ( .IN1(data1[11]), .IN2(n8), .IN3(data0[11]), .IN4(n7), .IN5(
        data2[11]), .IN6(n6), .Q(data_o[11]) );
  AO222X1 U18 ( .IN1(data1[10]), .IN2(n8), .IN3(data0[10]), .IN4(n7), .IN5(
        data2[10]), .IN6(n6), .Q(data_o[10]) );
  AO222X1 U19 ( .IN1(data1[0]), .IN2(n8), .IN3(data0[0]), .IN4(n7), .IN5(
        data2[0]), .IN6(n6), .Q(data_o[0]) );
  INVX0 U2 ( .INP(select0), .ZN(n2) );
  INVX0 U3 ( .INP(select1), .ZN(n1) );
  AND3X1 U20 ( .IN1(n2), .IN2(n1), .IN3(select2), .Q(n6) );
  NOR3X0 U21 ( .IN1(select1), .IN2(select2), .IN3(n2), .QN(n7) );
  NOR3X0 U22 ( .IN1(select0), .IN2(select2), .IN3(n1), .QN(n8) );
endmodule


module mux3_1_2 ( data0, data1, data2, select0, select1, select2, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  output [15:0] data_o;
  input select0, select1, select2;
  wire   n1, n2, n6, n7, n8;

  AO222X1 U4 ( .IN1(data1[9]), .IN2(n8), .IN3(data0[9]), .IN4(n7), .IN5(
        data2[9]), .IN6(n6), .Q(data_o[9]) );
  AO222X1 U5 ( .IN1(data1[8]), .IN2(n8), .IN3(data0[8]), .IN4(n7), .IN5(
        data2[8]), .IN6(n6), .Q(data_o[8]) );
  AO222X1 U6 ( .IN1(data1[7]), .IN2(n8), .IN3(data0[7]), .IN4(n7), .IN5(
        data2[7]), .IN6(n6), .Q(data_o[7]) );
  AO222X1 U7 ( .IN1(data1[6]), .IN2(n8), .IN3(data0[6]), .IN4(n7), .IN5(
        data2[6]), .IN6(n6), .Q(data_o[6]) );
  AO222X1 U8 ( .IN1(data1[5]), .IN2(n8), .IN3(data0[5]), .IN4(n7), .IN5(
        data2[5]), .IN6(n6), .Q(data_o[5]) );
  AO222X1 U9 ( .IN1(data1[4]), .IN2(n8), .IN3(data0[4]), .IN4(n7), .IN5(
        data2[4]), .IN6(n6), .Q(data_o[4]) );
  AO222X1 U10 ( .IN1(data1[3]), .IN2(n8), .IN3(data0[3]), .IN4(n7), .IN5(
        data2[3]), .IN6(n6), .Q(data_o[3]) );
  AO222X1 U11 ( .IN1(data1[2]), .IN2(n8), .IN3(data0[2]), .IN4(n7), .IN5(
        data2[2]), .IN6(n6), .Q(data_o[2]) );
  AO222X1 U12 ( .IN1(data1[1]), .IN2(n8), .IN3(data0[1]), .IN4(n7), .IN5(
        data2[1]), .IN6(n6), .Q(data_o[1]) );
  AO222X1 U13 ( .IN1(data1[15]), .IN2(n8), .IN3(data0[15]), .IN4(n7), .IN5(
        data2[15]), .IN6(n6), .Q(data_o[15]) );
  AO222X1 U14 ( .IN1(data1[14]), .IN2(n8), .IN3(data0[14]), .IN4(n7), .IN5(
        data2[14]), .IN6(n6), .Q(data_o[14]) );
  AO222X1 U15 ( .IN1(data1[13]), .IN2(n8), .IN3(data0[13]), .IN4(n7), .IN5(
        data2[13]), .IN6(n6), .Q(data_o[13]) );
  AO222X1 U16 ( .IN1(data1[12]), .IN2(n8), .IN3(data0[12]), .IN4(n7), .IN5(
        data2[12]), .IN6(n6), .Q(data_o[12]) );
  AO222X1 U17 ( .IN1(data1[11]), .IN2(n8), .IN3(data0[11]), .IN4(n7), .IN5(
        data2[11]), .IN6(n6), .Q(data_o[11]) );
  AO222X1 U18 ( .IN1(data1[10]), .IN2(n8), .IN3(data0[10]), .IN4(n7), .IN5(
        data2[10]), .IN6(n6), .Q(data_o[10]) );
  AO222X1 U19 ( .IN1(data1[0]), .IN2(n8), .IN3(data0[0]), .IN4(n7), .IN5(
        data2[0]), .IN6(n6), .Q(data_o[0]) );
  INVX0 U2 ( .INP(select0), .ZN(n2) );
  INVX0 U3 ( .INP(select1), .ZN(n1) );
  AND3X1 U20 ( .IN1(n2), .IN2(n1), .IN3(select2), .Q(n6) );
  NOR3X0 U21 ( .IN1(select1), .IN2(select2), .IN3(n2), .QN(n7) );
  NOR3X0 U22 ( .IN1(select0), .IN2(select2), .IN3(n1), .QN(n8) );
endmodule



    module node4_NODE_X3_NODE_Y1I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__I_node_2_node_interface__ ( 
        \clk.clk , \reset.reset , \local_node.clk , 
        \local_node.buffer_full_in , \local_node.buffer_full_out , 
        \local_node.receiving_data , \local_node.sending_data , 
        \local_node.data_in , \local_node.data_out , \node_0.clk , 
        \node_0.buffer_full_in , \node_0.buffer_full_out , 
        \node_0.receiving_data , \node_0.sending_data , \node_0.data_in , 
        \node_0.data_out , \node_1.clk , \node_1.buffer_full_in , 
        \node_1.buffer_full_out , \node_1.receiving_data , 
        \node_1.sending_data , \node_1.data_in , \node_1.data_out , 
        \node_2.clk , \node_2.buffer_full_in , \node_2.buffer_full_out , 
        \node_2.receiving_data , \node_2.sending_data , \node_2.data_in , 
        \node_2.data_out  );
  input [15:0] \local_node.data_in ;
  output [15:0] \local_node.data_out ;
  input [15:0] \node_0.data_in ;
  output [15:0] \node_0.data_out ;
  input [15:0] \node_1.data_in ;
  output [15:0] \node_1.data_out ;
  input [15:0] \node_2.data_in ;
  output [15:0] \node_2.data_out ;
  input \clk.clk , \reset.reset , \local_node.buffer_full_in ,
         \local_node.receiving_data , \node_0.buffer_full_in ,
         \node_0.receiving_data , \node_1.buffer_full_in ,
         \node_1.receiving_data , \node_2.buffer_full_in ,
         \node_2.receiving_data ;
  output \local_node.buffer_full_out , \local_node.sending_data ,
         \node_0.buffer_full_out , \node_0.sending_data ,
         \node_1.buffer_full_out , \node_1.sending_data ,
         \node_2.buffer_full_out , \node_2.sending_data ;
  inout \local_node.clk ,  \node_0.clk ,  \node_1.clk ,  \node_2.clk ;
  wire   \buffer_out[3][15] , \buffer_out[3][14] , \buffer_out[3][13] ,
         \buffer_out[3][12] , \buffer_out[3][11] , \buffer_out[3][10] ,
         \buffer_out[3][9] , \buffer_out[3][8] , \buffer_out[3][7] ,
         \buffer_out[3][6] , \buffer_out[3][5] , \buffer_out[3][4] ,
         \buffer_out[3][3] , \buffer_out[3][2] , \buffer_out[3][1] ,
         \buffer_out[3][0] , \buffer_out[2][15] , \buffer_out[2][14] ,
         \buffer_out[2][13] , \buffer_out[2][12] , \buffer_out[2][11] ,
         \buffer_out[2][10] , \buffer_out[2][9] , \buffer_out[2][8] ,
         \buffer_out[2][7] , \buffer_out[2][6] , \buffer_out[2][5] ,
         \buffer_out[2][4] , \buffer_out[2][3] , \buffer_out[2][2] ,
         \buffer_out[2][1] , \buffer_out[2][0] , \buffer_out[1][15] ,
         \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] ,
         \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] ,
         \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] ,
         \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] ,
         \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] ,
         \buffer_out[0][15] , \buffer_out[0][14] , \buffer_out[0][13] ,
         \buffer_out[0][12] , \buffer_out[0][11] , \buffer_out[0][10] ,
         \buffer_out[0][9] , \buffer_out[0][8] , \buffer_out[0][7] ,
         \buffer_out[0][6] , \buffer_out[0][5] , \buffer_out[0][4] ,
         \buffer_out[0][3] , \buffer_out[0][2] , \buffer_out[0][1] ,
         \buffer_out[0][0] , \next_buffer_out[3][15] ,
         \next_buffer_out[3][14] , \next_buffer_out[3][13] ,
         \next_buffer_out[3][12] , \next_buffer_out[3][11] ,
         \next_buffer_out[3][10] , \next_buffer_out[3][9] ,
         \next_buffer_out[3][8] , \next_buffer_out[3][7] ,
         \next_buffer_out[3][6] , \next_buffer_out[3][5] ,
         \next_buffer_out[3][4] , \next_buffer_out[3][3] ,
         \next_buffer_out[3][2] , \next_buffer_out[3][1] ,
         \next_buffer_out[3][0] , \next_buffer_out[2][15] ,
         \next_buffer_out[2][14] , \next_buffer_out[2][13] ,
         \next_buffer_out[2][12] , \next_buffer_out[2][11] ,
         \next_buffer_out[2][10] , \next_buffer_out[2][9] ,
         \next_buffer_out[2][8] , \next_buffer_out[2][7] ,
         \next_buffer_out[2][6] , \next_buffer_out[2][5] ,
         \next_buffer_out[2][4] , \next_buffer_out[2][3] ,
         \next_buffer_out[2][2] , \next_buffer_out[2][1] ,
         \next_buffer_out[2][0] , \next_buffer_out[1][15] ,
         \next_buffer_out[1][14] , \next_buffer_out[1][13] ,
         \next_buffer_out[1][12] , \next_buffer_out[1][11] ,
         \next_buffer_out[1][10] , \next_buffer_out[1][9] ,
         \next_buffer_out[1][8] , \next_buffer_out[1][7] ,
         \next_buffer_out[1][6] , \next_buffer_out[1][5] ,
         \next_buffer_out[1][4] , \next_buffer_out[1][3] ,
         \next_buffer_out[1][2] , \next_buffer_out[1][1] ,
         \next_buffer_out[1][0] , \next_buffer_out[0][15] ,
         \next_buffer_out[0][14] , \next_buffer_out[0][13] ,
         \next_buffer_out[0][12] , \next_buffer_out[0][11] ,
         \next_buffer_out[0][10] , \next_buffer_out[0][9] ,
         \next_buffer_out[0][8] , \next_buffer_out[0][7] ,
         \next_buffer_out[0][6] , \next_buffer_out[0][5] ,
         \next_buffer_out[0][4] , \next_buffer_out[0][3] ,
         \next_buffer_out[0][2] , \next_buffer_out[0][1] ,
         \next_buffer_out[0][0] ;
  wire   [3:0] buffer_full_in;
  wire   [3:0] receiving_data;
  wire   [3:0] pop_v;
  wire   [3:0] data_valid;
  wire   [3:0] next_data_valid;
  wire   [1:0] grant_0;
  wire   [1:0] grant_1;
  wire   [2:0] grant_2;
  wire   [2:0] grant_3;
  tri   \local_node.buffer_full_in ;
  tri   \local_node.buffer_full_out ;
  tri   \local_node.receiving_data ;
  tri   \local_node.sending_data ;
  tri   [15:0] \local_node.data_in ;
  tri   [15:0] \local_node.data_out ;

  converter_out_I_n_node_interface_dut_ c3 ( .\n.buffer_full_in (
        \local_node.buffer_full_in ), .\n.receiving_data (
        \local_node.receiving_data ), .\n.data_in (\local_node.data_in ), 
        .\n.buffer_full_out (\local_node.buffer_full_out ), .\n.sending_data (
        \local_node.sending_data ), .\n.data_out (\local_node.data_out ), 
        .buffer_full_in(1'b0), .receiving_data(1'b0), .data_in({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  fifo_kev_27 \genblk1[0].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[0]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[0]), .data_out({\buffer_out[0][15] , 
        \buffer_out[0][14] , \buffer_out[0][13] , \buffer_out[0][12] , 
        \buffer_out[0][11] , \buffer_out[0][10] , \buffer_out[0][9] , 
        \buffer_out[0][8] , \buffer_out[0][7] , \buffer_out[0][6] , 
        \buffer_out[0][5] , \buffer_out[0][4] , \buffer_out[0][3] , 
        \buffer_out[0][2] , \buffer_out[0][1] , \buffer_out[0][0] }), 
        .next_data_out({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] , 
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .next_data_valid(
        next_data_valid[0]) );
  address_counter_27 \genblk1[0].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] }), 
        .buffer_data_valid(next_data_valid[0]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .buffer_pop(
        pop_v[0]), .receiving_data(1'b0) );
  fifo_kev_26 \genblk1[1].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[1]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[1]), .data_out({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), 
        .next_data_out({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] , 
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .next_data_valid(
        next_data_valid[1]) );
  address_counter_26 \genblk1[1].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] }), 
        .buffer_data_valid(next_data_valid[1]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .buffer_pop(
        pop_v[1]), .receiving_data(1'b0) );
  fifo_kev_25 \genblk1[2].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[2]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[2]), .data_out({\buffer_out[2][15] , 
        \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] , 
        \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] , 
        \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] , 
        \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] , 
        \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] }), 
        .next_data_out({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] , 
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .next_data_valid(
        next_data_valid[2]) );
  address_counter_25 \genblk1[2].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] }), 
        .buffer_data_valid(next_data_valid[2]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .buffer_pop(
        pop_v[2]), .receiving_data(1'b0) );
  fifo_kev_24 \genblk1[3].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[3]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[3]), .data_out({\buffer_out[3][15] , 
        \buffer_out[3][14] , \buffer_out[3][13] , \buffer_out[3][12] , 
        \buffer_out[3][11] , \buffer_out[3][10] , \buffer_out[3][9] , 
        \buffer_out[3][8] , \buffer_out[3][7] , \buffer_out[3][6] , 
        \buffer_out[3][5] , \buffer_out[3][4] , \buffer_out[3][3] , 
        \buffer_out[3][2] , \buffer_out[3][1] , \buffer_out[3][0] }), 
        .next_data_out({\next_buffer_out[3][15] , \next_buffer_out[3][14] , 
        \next_buffer_out[3][13] , \next_buffer_out[3][12] , 
        \next_buffer_out[3][11] , \next_buffer_out[3][10] , 
        \next_buffer_out[3][9] , \next_buffer_out[3][8] , 
        \next_buffer_out[3][7] , \next_buffer_out[3][6] , 
        \next_buffer_out[3][5] , \next_buffer_out[3][4] , 
        \next_buffer_out[3][3] , \next_buffer_out[3][2] , 
        \next_buffer_out[3][1] , \next_buffer_out[3][0] }), .next_data_valid(
        next_data_valid[3]) );
  address_counter_24 \genblk1[3].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[3][15] , \next_buffer_out[3][14] , 
        \next_buffer_out[3][13] , \next_buffer_out[3][12] , 
        \next_buffer_out[3][11] , \next_buffer_out[3][10] , 
        \next_buffer_out[3][9] , \next_buffer_out[3][8] }), 
        .buffer_data_valid(next_data_valid[3]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[3][7] , \next_buffer_out[3][6] , 
        \next_buffer_out[3][5] , \next_buffer_out[3][4] , 
        \next_buffer_out[3][3] , \next_buffer_out[3][2] , 
        \next_buffer_out[3][1] , \next_buffer_out[3][0] }), .buffer_pop(
        pop_v[3]), .receiving_data(1'b0) );
  converter_in_I_n_node_interface_dut__9 \genblk2.c0  ( .\n.buffer_full_in (
        \node_0.buffer_full_in ), .\n.receiving_data (\node_0.receiving_data ), 
        .\n.data_in (\node_0.data_in ), .\n.buffer_full_out (
        \node_0.buffer_full_out ), .\n.sending_data (\node_0.sending_data ), 
        .\n.data_out (\node_0.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_out_I_n_node_interface_dut_ \genblk2.c1  ( .\n.buffer_full_in (
        \node_1.buffer_full_in ), .\n.receiving_data (\node_1.receiving_data ), 
        .\n.data_in (\node_1.data_in ), .\n.buffer_full_out (
        \node_1.buffer_full_out ), .\n.sending_data (\node_1.sending_data ), 
        .\n.data_out (\node_1.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_out_I_n_node_interface_dut_ \genblk2.c2  ( .\n.buffer_full_in (
        \node_2.buffer_full_in ), .\n.receiving_data (\node_2.receiving_data ), 
        .\n.data_in (\node_2.data_in ), .\n.buffer_full_out (
        \node_2.buffer_full_out ), .\n.sending_data (\node_2.sending_data ), 
        .\n.data_out (\node_2.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  controller4_edge_e_1 \genblk2.e  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .packet_addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .local_addr({1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1}), 
        .packet_valid(data_valid), .buffer_full_in({1'b0, 1'b0, 1'b0, 1'b0}), 
        .grant_0(grant_0), .grant_1(grant_1), .grant_2(grant_2), .grant_3(
        grant_3), .pop_v(pop_v) );
  mux2_1_11 \genblk2.mux_n  ( .data0({\buffer_out[1][15] , \buffer_out[1][14] , 
        \buffer_out[1][13] , \buffer_out[1][12] , \buffer_out[1][11] , 
        \buffer_out[1][10] , \buffer_out[1][9] , \buffer_out[1][8] , 
        \buffer_out[1][7] , \buffer_out[1][6] , \buffer_out[1][5] , 
        \buffer_out[1][4] , \buffer_out[1][3] , \buffer_out[1][2] , 
        \buffer_out[1][1] , \buffer_out[1][0] }), .data1({\buffer_out[3][15] , 
        \buffer_out[3][14] , \buffer_out[3][13] , \buffer_out[3][12] , 
        \buffer_out[3][11] , \buffer_out[3][10] , \buffer_out[3][9] , 
        \buffer_out[3][8] , \buffer_out[3][7] , \buffer_out[3][6] , 
        \buffer_out[3][5] , \buffer_out[3][4] , \buffer_out[3][3] , 
        \buffer_out[3][2] , \buffer_out[3][1] , \buffer_out[3][0] }), 
        .select0(grant_0[0]), .select1(grant_0[1]) );
  mux2_1_10 \genblk2.mux_s  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[3][15] , 
        \buffer_out[3][14] , \buffer_out[3][13] , \buffer_out[3][12] , 
        \buffer_out[3][11] , \buffer_out[3][10] , \buffer_out[3][9] , 
        \buffer_out[3][8] , \buffer_out[3][7] , \buffer_out[3][6] , 
        \buffer_out[3][5] , \buffer_out[3][4] , \buffer_out[3][3] , 
        \buffer_out[3][2] , \buffer_out[3][1] , \buffer_out[3][0] }), 
        .select0(grant_1[0]), .select1(grant_1[1]) );
  mux3_1_3 \genblk2.mux_w  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[3][15] , \buffer_out[3][14] , \buffer_out[3][13] , 
        \buffer_out[3][12] , \buffer_out[3][11] , \buffer_out[3][10] , 
        \buffer_out[3][9] , \buffer_out[3][8] , \buffer_out[3][7] , 
        \buffer_out[3][6] , \buffer_out[3][5] , \buffer_out[3][4] , 
        \buffer_out[3][3] , \buffer_out[3][2] , \buffer_out[3][1] , 
        \buffer_out[3][0] }), .select0(grant_2[0]), .select1(grant_2[1]), 
        .select2(grant_2[2]) );
  mux3_1_2 \genblk2.mux_l  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[2][15] , \buffer_out[2][14] , \buffer_out[2][13] , 
        \buffer_out[2][12] , \buffer_out[2][11] , \buffer_out[2][10] , 
        \buffer_out[2][9] , \buffer_out[2][8] , \buffer_out[2][7] , 
        \buffer_out[2][6] , \buffer_out[2][5] , \buffer_out[2][4] , 
        \buffer_out[2][3] , \buffer_out[2][2] , \buffer_out[2][1] , 
        \buffer_out[2][0] }), .select0(grant_3[0]), .select1(grant_3[1]), 
        .select2(grant_3[2]) );
endmodule


module fifo_kev_23 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_47 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_23 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_47 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_46 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_23 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_46 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_23_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_23 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_23 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_23 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_23_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_22 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_45 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_22 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_45 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_44 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_22 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_44 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_22_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_22 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_22 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_22 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_22_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_21 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_43 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_21 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_43 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_42 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_21 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_42 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_21_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_21 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_21 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_21 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_21_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_20 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_41 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_20 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_41 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_40 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_20 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_40 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_20_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_20 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_20 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_20 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_20_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module converter_in_I_n_node_interface_dut__8 ( \n.buffer_full_in , 
        \n.receiving_data , \n.data_in , \n.buffer_full_out , \n.sending_data , 
        \n.data_out , buffer_full_out, sending_data, data_out, buffer_full_in, 
        receiving_data, data_in );
  input [15:0] \n.data_in ;
  output [15:0] \n.data_out ;
  output [15:0] data_out;
  input [15:0] data_in;
  input \n.buffer_full_in , \n.receiving_data , buffer_full_in, receiving_data;
  output \n.buffer_full_out , \n.sending_data , buffer_full_out, sending_data;
  wire   \n.buffer_full_in , \n.receiving_data , buffer_full_in,
         receiving_data;
  assign buffer_full_out = \n.buffer_full_in ;
  assign sending_data = \n.receiving_data ;
  assign data_out[15] = \n.data_in  [15];
  assign data_out[14] = \n.data_in  [14];
  assign data_out[13] = \n.data_in  [13];
  assign data_out[12] = \n.data_in  [12];
  assign data_out[11] = \n.data_in  [11];
  assign data_out[10] = \n.data_in  [10];
  assign data_out[9] = \n.data_in  [9];
  assign data_out[8] = \n.data_in  [8];
  assign data_out[7] = \n.data_in  [7];
  assign data_out[6] = \n.data_in  [6];
  assign data_out[5] = \n.data_in  [5];
  assign data_out[4] = \n.data_in  [4];
  assign data_out[3] = \n.data_in  [3];
  assign data_out[2] = \n.data_in  [2];
  assign data_out[1] = \n.data_in  [1];
  assign data_out[0] = \n.data_in  [0];
  assign \n.buffer_full_out  = buffer_full_in;
  assign \n.sending_data  = receiving_data;
  assign \n.data_out  [15] = data_in[15];
  assign \n.data_out  [14] = data_in[14];
  assign \n.data_out  [13] = data_in[13];
  assign \n.data_out  [12] = data_in[12];
  assign \n.data_out  [11] = data_in[11];
  assign \n.data_out  [10] = data_in[10];
  assign \n.data_out  [9] = data_in[9];
  assign \n.data_out  [8] = data_in[8];
  assign \n.data_out  [7] = data_in[7];
  assign \n.data_out  [6] = data_in[6];
  assign \n.data_out  [5] = data_in[5];
  assign \n.data_out  [4] = data_in[4];
  assign \n.data_out  [3] = data_in[3];
  assign \n.data_out  [2] = data_in[2];
  assign \n.data_out  [1] = data_in[1];
  assign \n.data_out  [0] = data_in[0];

endmodule


module flipflop_BITS2_9 ( clk, data_i, data_o );
  input [1:0] data_i;
  output [1:0] data_o;
  input clk;


  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS2_9 ( clk, enable_i, reset, data_i, data_o );
  input [1:0] data_i;
  input [1:0] data_o;
  input clk, enable_i, reset;
  wire   n10, n11, n1, n5, n7, n8, n9;
  wire   [1:0] write_data;

  AOI22X1 U5 ( .IN1(enable_i), .IN2(data_i[1]), .IN3(n10), .IN4(n1), .QN(n9)
         );
  AOI22X1 U6 ( .IN1(data_i[0]), .IN2(enable_i), .IN3(n11), .IN4(n1), .QN(n8)
         );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n9), .QN(write_data[1]) );
  NOR2X0 U4 ( .IN1(reset), .IN2(n8), .QN(write_data[0]) );
  AND2X1 U7 ( .IN1(data_o[1]), .IN2(n7), .Q(n10) );
  AND2X1 U8 ( .IN1(data_o[0]), .IN2(n5), .Q(n11) );
  flipflop_BITS2_9 FF ( .clk(clk), .data_i(write_data), .data_o({n7, n5}) );
endmodule


module flipflop_BITS1_37 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_37 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_37 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter2_9 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [1:0] request;
  output [1:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   tail_en, n1, n2;
  wire   [1:0] req_i;
  wire   [1:0] req_o;

  AND3X1 U10 ( .IN1(request[1]), .IN2(n1), .IN3(n2), .Q(grant[1]) );
  AND3X1 U11 ( .IN1(request[0]), .IN2(n2), .IN3(request[1]), .Q(tail_en) );
  INVX0 U6 ( .INP(request[0]), .ZN(n1) );
  NOR2X0 U7 ( .IN1(buffer_full_i), .IN2(n1), .QN(grant[0]) );
  INVX0 U8 ( .INP(buffer_full_i), .ZN(n2) );
  OA21X1 U9 ( .IN1(request[1]), .IN2(request[0]), .IN3(n2), .Q(grant_v_o) );
  register_BITS2_9 req_record ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i({1'b1, 1'b0}), .data_o({1'b0, 1'b0}) );
  register_BITS1_37 tail ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i(1'b1), .data_o(1'b0) );
endmodule


module flipflop_BITS2_8 ( clk, data_i, data_o );
  input [1:0] data_i;
  output [1:0] data_o;
  input clk;


  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS2_8 ( clk, enable_i, reset, data_i, data_o );
  input [1:0] data_i;
  input [1:0] data_o;
  input clk, enable_i, reset;
  wire   n10, n11, n1, n5, n7, n8, n9;
  wire   [1:0] write_data;

  AOI22X1 U5 ( .IN1(enable_i), .IN2(data_i[1]), .IN3(n10), .IN4(n1), .QN(n9)
         );
  AOI22X1 U6 ( .IN1(data_i[0]), .IN2(enable_i), .IN3(n11), .IN4(n1), .QN(n8)
         );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n9), .QN(write_data[1]) );
  NOR2X0 U4 ( .IN1(reset), .IN2(n8), .QN(write_data[0]) );
  AND2X1 U7 ( .IN1(data_o[1]), .IN2(n7), .Q(n10) );
  AND2X1 U8 ( .IN1(data_o[0]), .IN2(n5), .Q(n11) );
  flipflop_BITS2_8 FF ( .clk(clk), .data_i(write_data), .data_o({n7, n5}) );
endmodule


module flipflop_BITS1_36 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_36 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_36 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter2_8 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [1:0] request;
  output [1:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   tail_en, n1, n2;
  wire   [1:0] req_i;
  wire   [1:0] req_o;

  AND3X1 U10 ( .IN1(request[1]), .IN2(n1), .IN3(n2), .Q(grant[1]) );
  AND3X1 U11 ( .IN1(request[0]), .IN2(n2), .IN3(request[1]), .Q(tail_en) );
  INVX0 U6 ( .INP(request[0]), .ZN(n1) );
  NOR2X0 U7 ( .IN1(buffer_full_i), .IN2(n1), .QN(grant[0]) );
  INVX0 U8 ( .INP(buffer_full_i), .ZN(n2) );
  OA21X1 U9 ( .IN1(request[1]), .IN2(request[0]), .IN3(n2), .Q(grant_v_o) );
  register_BITS2_8 req_record ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i({1'b1, 1'b0}), .data_o({1'b0, 1'b0}) );
  register_BITS1_36 tail ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i(1'b1), .data_o(1'b0) );
endmodule


module flipflop_BITS3_3 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_3 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_3 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS3_2 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_2 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_2 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS1_35 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_35 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_35 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_34 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_34 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_34 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter3_1 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [2:0] request;
  output [2:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[1][2] , \req_i[1][1] , \req_i[1][0] , \req_i[0][2] ,
         \req_i[0][1] , tail_en, N99, N100, N101, N110, N111, N118, N119, N120,
         N121, n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [1:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N99 = request[0];
  assign N100 = request[1];
  assign N101 = request[2];

  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(N111), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(N110), .Q(\req_i[0][1] ) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N121), .D(tail_en), .Q(req_en[0]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N120), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N119), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N118), .Q(grant[0]) );
  AND2X1 U20 ( .IN1(n8), .IN2(N101), .Q(n7) );
  OR3X1 U21 ( .IN1(n3), .IN2(N111), .IN3(n6), .Q(N121) );
  NOR3X0 U22 ( .IN1(N99), .IN2(N100), .IN3(n6), .QN(N120) );
  NOR3X0 U23 ( .IN1(n2), .IN2(N99), .IN3(n6), .QN(N119) );
  NAND3X0 U24 ( .IN1(n2), .IN2(n3), .IN3(n1), .QN(n5) );
  AO22X1 U25 ( .IN1(N100), .IN2(N101), .IN3(N99), .IN4(N101), .Q(N111) );
  INVX0 U10 ( .INP(N101), .ZN(n3) );
  NAND2X1 U11 ( .IN1(n5), .IN2(n4), .QN(n6) );
  INVX0 U12 ( .INP(N99), .ZN(n1) );
  INVX0 U13 ( .INP(N100), .ZN(n2) );
  INVX0 U14 ( .INP(buffer_full_i), .ZN(n4) );
  NAND2X1 U15 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NOR2X0 U16 ( .IN1(n1), .IN2(n6), .QN(N118) );
  NOR2X0 U17 ( .IN1(n1), .IN2(n2), .QN(N110) );
  OA21X1 U18 ( .IN1(N110), .IN2(n7), .IN3(n4), .Q(tail_en) );
  OA21X1 U19 ( .IN1(N101), .IN2(n8), .IN3(n4), .Q(grant_v_o) );
  register_BITS3_3 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][2] , \req_i[0][1] , 1'b0}), .data_o({
        1'b0, 1'b0, 1'b0}) );
  register_BITS3_2 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][2] , \req_i[1][1] , \req_i[1][0] }), 
        .data_o({1'b0, 1'b0, 1'b0}) );
  register_BITS1_35 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b1), .data_o(1'b0) );
  register_BITS1_34 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module flipflop_BITS3_1 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_1 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_1 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS3_0 ( clk, data_i, data_o );
  input [2:0] data_i;
  output [2:0] data_o;
  input clk;


  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS3_0 ( clk, enable_i, reset, data_i, data_o );
  input [2:0] data_i;
  input [2:0] data_o;
  input clk, enable_i, reset;
  wire   n12, n13, n14, n1, n5, n7, n9, n10, n11;
  wire   [2:0] write_data;

  AO22X1 U5 ( .IN1(data_i[2]), .IN2(n11), .IN3(n12), .IN4(n10), .Q(
        write_data[2]) );
  AO22X1 U6 ( .IN1(data_i[1]), .IN2(n11), .IN3(n13), .IN4(n10), .Q(
        write_data[1]) );
  AO22X1 U7 ( .IN1(data_i[0]), .IN2(n11), .IN3(n14), .IN4(n10), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n10) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n11) );
  AND2X1 U8 ( .IN1(data_o[2]), .IN2(n9), .Q(n12) );
  AND2X1 U9 ( .IN1(data_o[1]), .IN2(n7), .Q(n13) );
  AND2X1 U10 ( .IN1(data_o[0]), .IN2(n5), .Q(n14) );
  flipflop_BITS3_0 FF ( .clk(clk), .data_i(write_data), .data_o({n9, n7, n5})
         );
endmodule


module flipflop_BITS1_33 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_33 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_33 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_32 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_32 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_32 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter3_0 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [2:0] request;
  output [2:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[1][2] , \req_i[1][1] , \req_i[1][0] , \req_i[0][2] ,
         \req_i[0][1] , tail_en, N99, N100, N101, N110, N111, N118, N119, N120,
         N121, n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [1:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N99 = request[0];
  assign N100 = request[1];
  assign N101 = request[2];

  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(N111), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(N110), .Q(\req_i[0][1] ) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N121), .D(tail_en), .Q(req_en[0]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N120), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N119), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N118), .Q(grant[0]) );
  AND2X1 U20 ( .IN1(n8), .IN2(N101), .Q(n7) );
  OR3X1 U21 ( .IN1(n3), .IN2(N111), .IN3(n6), .Q(N121) );
  NOR3X0 U22 ( .IN1(N99), .IN2(N100), .IN3(n6), .QN(N120) );
  NOR3X0 U23 ( .IN1(n2), .IN2(N99), .IN3(n6), .QN(N119) );
  NAND3X0 U24 ( .IN1(n2), .IN2(n3), .IN3(n1), .QN(n5) );
  AO22X1 U25 ( .IN1(N100), .IN2(N101), .IN3(N99), .IN4(N101), .Q(N111) );
  INVX0 U10 ( .INP(N101), .ZN(n3) );
  NAND2X1 U11 ( .IN1(n5), .IN2(n4), .QN(n6) );
  INVX0 U12 ( .INP(N99), .ZN(n1) );
  INVX0 U13 ( .INP(N100), .ZN(n2) );
  INVX0 U14 ( .INP(buffer_full_i), .ZN(n4) );
  NAND2X1 U15 ( .IN1(n1), .IN2(n2), .QN(n8) );
  NOR2X0 U16 ( .IN1(n1), .IN2(n6), .QN(N118) );
  NOR2X0 U17 ( .IN1(n1), .IN2(n2), .QN(N110) );
  OA21X1 U18 ( .IN1(N110), .IN2(n7), .IN3(n4), .Q(tail_en) );
  OA21X1 U19 ( .IN1(N101), .IN2(n8), .IN3(n4), .Q(grant_v_o) );
  register_BITS3_1 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][2] , \req_i[0][1] , 1'b0}), .data_o({
        1'b0, 1'b0, 1'b0}) );
  register_BITS3_0 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][2] , \req_i[1][1] , \req_i[1][0] }), 
        .data_o({1'b0, 1'b0, 1'b0}) );
  register_BITS1_33 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b1), .data_o(1'b0) );
  register_BITS1_32 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module dccl_23 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_22 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_21 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_20 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module controller4_edge_e_0 ( clk, rst, .packet_addr({\packet_addr[3][7] , 
        \packet_addr[3][6] , \packet_addr[3][5] , \packet_addr[3][4] , 
        \packet_addr[3][3] , \packet_addr[3][2] , \packet_addr[3][1] , 
        \packet_addr[3][0] , \packet_addr[2][7] , \packet_addr[2][6] , 
        \packet_addr[2][5] , \packet_addr[2][4] , \packet_addr[2][3] , 
        \packet_addr[2][2] , \packet_addr[2][1] , \packet_addr[2][0] , 
        \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] , 
        \packet_addr[1][4] , \packet_addr[1][3] , \packet_addr[1][2] , 
        \packet_addr[1][1] , \packet_addr[1][0] , \packet_addr[0][7] , 
        \packet_addr[0][6] , \packet_addr[0][5] , \packet_addr[0][4] , 
        \packet_addr[0][3] , \packet_addr[0][2] , \packet_addr[0][1] , 
        \packet_addr[0][0] }), local_addr, packet_valid, buffer_full_in, 
        grant_0, grant_1, grant_2, grant_3, grant_v, pop_v );
  input [7:0] local_addr;
  input [3:0] packet_valid;
  input [3:0] buffer_full_in;
  output [1:0] grant_0;
  output [1:0] grant_1;
  output [2:0] grant_2;
  output [2:0] grant_3;
  output [3:0] grant_v;
  output [3:0] pop_v;
  input clk, rst, \packet_addr[3][7] , \packet_addr[3][6] ,
         \packet_addr[3][5] , \packet_addr[3][4] , \packet_addr[3][3] ,
         \packet_addr[3][2] , \packet_addr[3][1] , \packet_addr[3][0] ,
         \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] ,
         \packet_addr[2][4] , \packet_addr[2][3] , \packet_addr[2][2] ,
         \packet_addr[2][1] , \packet_addr[2][0] , \packet_addr[1][7] ,
         \packet_addr[1][6] , \packet_addr[1][5] , \packet_addr[1][4] ,
         \packet_addr[1][3] , \packet_addr[1][2] , \packet_addr[1][1] ,
         \packet_addr[1][0] , \packet_addr[0][7] , \packet_addr[0][6] ,
         \packet_addr[0][5] , \packet_addr[0][4] , \packet_addr[0][3] ,
         \packet_addr[0][2] , \packet_addr[0][1] , \packet_addr[0][0] ;
  wire   \grant_3[2] , \request[3][2] , \request[3][1] , \request[3][0] ,
         \request[2][2] , \request[2][1] , \request[2][0] , \request[1][1] ,
         \request[1][0] , \request[0][1] , \request[0][0] ;
  assign pop_v[2] = \grant_3[2] ;
  assign grant_3[2] = \grant_3[2] ;

  OR3X1 U1 ( .IN1(grant_2[2]), .IN2(grant_1[1]), .IN3(grant_0[1]), .Q(pop_v[3]) );
  OR3X1 U2 ( .IN1(grant_3[1]), .IN2(grant_2[1]), .IN3(grant_0[0]), .Q(pop_v[1]) );
  OR3X1 U3 ( .IN1(grant_3[0]), .IN2(grant_2[0]), .IN3(grant_1[0]), .Q(pop_v[0]) );
  arbiter2_9 arbiter_n ( .clk(clk), .rst(rst), .request({\request[0][1] , 
        \request[0][0] }), .buffer_full_i(buffer_full_in[0]), .grant(grant_0), 
        .grant_v_o(grant_v[0]) );
  arbiter2_8 arbiter_s ( .clk(clk), .rst(rst), .request({\request[1][1] , 
        \request[1][0] }), .buffer_full_i(buffer_full_in[1]), .grant(grant_1), 
        .grant_v_o(grant_v[1]) );
  arbiter3_1 arbiter_w ( .clk(clk), .rst(rst), .request({\request[2][2] , 
        \request[2][1] , \request[2][0] }), .buffer_full_i(buffer_full_in[2]), 
        .grant(grant_2), .grant_v_o(grant_v[2]) );
  arbiter3_0 arbiter_l ( .clk(clk), .rst(rst), .request({\request[3][2] , 
        \request[3][1] , \request[3][0] }), .buffer_full_i(buffer_full_in[3]), 
        .grant({\grant_3[2] , grant_3[1:0]}), .grant_v_o(grant_v[3]) );
  dccl_23 dccl_n ( .packet_addr_y_i({\packet_addr[0][3] , \packet_addr[0][2] , 
        \packet_addr[0][1] , \packet_addr[0][0] }), .packet_addr_x_i({
        \packet_addr[0][7] , \packet_addr[0][6] , \packet_addr[0][5] , 
        \packet_addr[0][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[0]), 
        .south_req(\request[1][0] ), .west_req(\request[2][0] ), .local_req(
        \request[3][0] ) );
  dccl_22 dccl_s ( .packet_addr_y_i({\packet_addr[1][3] , \packet_addr[1][2] , 
        \packet_addr[1][1] , \packet_addr[1][0] }), .packet_addr_x_i({
        \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] , 
        \packet_addr[1][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[1]), 
        .north_req(\request[0][0] ), .west_req(\request[2][1] ), .local_req(
        \request[3][1] ) );
  dccl_21 dccl_w ( .packet_addr_y_i({\packet_addr[2][3] , \packet_addr[2][2] , 
        \packet_addr[2][1] , \packet_addr[2][0] }), .packet_addr_x_i({
        \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] , 
        \packet_addr[2][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[2]), 
        .local_req(\request[3][2] ) );
  dccl_20 dccl_l ( .packet_addr_y_i({\packet_addr[3][3] , \packet_addr[3][2] , 
        \packet_addr[3][1] , \packet_addr[3][0] }), .packet_addr_x_i({
        \packet_addr[3][7] , \packet_addr[3][6] , \packet_addr[3][5] , 
        \packet_addr[3][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[3]), 
        .north_req(\request[0][1] ), .south_req(\request[1][1] ), .west_req(
        \request[2][2] ) );
endmodule


module mux2_1_9 ( data0, data1, select0, select1, data_o );
  input [15:0] data0;
  input [15:0] data1;
  output [15:0] data_o;
  input select0, select1;
  wire   n1, n4, n5;

  AO22X1 U4 ( .IN1(data1[9]), .IN2(n5), .IN3(data0[9]), .IN4(n4), .Q(data_o[9]) );
  AO22X1 U5 ( .IN1(data1[8]), .IN2(n5), .IN3(data0[8]), .IN4(n4), .Q(data_o[8]) );
  AO22X1 U6 ( .IN1(data1[7]), .IN2(n5), .IN3(data0[7]), .IN4(n4), .Q(data_o[7]) );
  AO22X1 U7 ( .IN1(data1[6]), .IN2(n5), .IN3(data0[6]), .IN4(n4), .Q(data_o[6]) );
  AO22X1 U8 ( .IN1(data1[5]), .IN2(n5), .IN3(data0[5]), .IN4(n4), .Q(data_o[5]) );
  AO22X1 U9 ( .IN1(data1[4]), .IN2(n5), .IN3(data0[4]), .IN4(n4), .Q(data_o[4]) );
  AO22X1 U10 ( .IN1(data1[3]), .IN2(n5), .IN3(data0[3]), .IN4(n4), .Q(
        data_o[3]) );
  AO22X1 U11 ( .IN1(data1[2]), .IN2(n5), .IN3(data0[2]), .IN4(n4), .Q(
        data_o[2]) );
  AO22X1 U12 ( .IN1(data1[1]), .IN2(n5), .IN3(data0[1]), .IN4(n4), .Q(
        data_o[1]) );
  AO22X1 U13 ( .IN1(data1[15]), .IN2(n5), .IN3(data0[15]), .IN4(n4), .Q(
        data_o[15]) );
  AO22X1 U14 ( .IN1(data1[14]), .IN2(n5), .IN3(data0[14]), .IN4(n4), .Q(
        data_o[14]) );
  AO22X1 U15 ( .IN1(data1[13]), .IN2(n5), .IN3(data0[13]), .IN4(n4), .Q(
        data_o[13]) );
  AO22X1 U16 ( .IN1(data1[12]), .IN2(n5), .IN3(data0[12]), .IN4(n4), .Q(
        data_o[12]) );
  AO22X1 U17 ( .IN1(data1[11]), .IN2(n5), .IN3(data0[11]), .IN4(n4), .Q(
        data_o[11]) );
  AO22X1 U18 ( .IN1(data1[10]), .IN2(n5), .IN3(data0[10]), .IN4(n4), .Q(
        data_o[10]) );
  AO22X1 U19 ( .IN1(data1[0]), .IN2(n5), .IN3(data0[0]), .IN4(n4), .Q(
        data_o[0]) );
  INVX0 U2 ( .INP(select1), .ZN(n1) );
  AND2X1 U3 ( .IN1(select0), .IN2(n1), .Q(n4) );
  NOR2X0 U20 ( .IN1(n1), .IN2(select0), .QN(n5) );
endmodule


module mux2_1_8 ( data0, data1, select0, select1, data_o );
  input [15:0] data0;
  input [15:0] data1;
  output [15:0] data_o;
  input select0, select1;
  wire   n1, n4, n5;

  AO22X1 U4 ( .IN1(data1[9]), .IN2(n5), .IN3(data0[9]), .IN4(n4), .Q(data_o[9]) );
  AO22X1 U5 ( .IN1(data1[8]), .IN2(n5), .IN3(data0[8]), .IN4(n4), .Q(data_o[8]) );
  AO22X1 U6 ( .IN1(data1[7]), .IN2(n5), .IN3(data0[7]), .IN4(n4), .Q(data_o[7]) );
  AO22X1 U7 ( .IN1(data1[6]), .IN2(n5), .IN3(data0[6]), .IN4(n4), .Q(data_o[6]) );
  AO22X1 U8 ( .IN1(data1[5]), .IN2(n5), .IN3(data0[5]), .IN4(n4), .Q(data_o[5]) );
  AO22X1 U9 ( .IN1(data1[4]), .IN2(n5), .IN3(data0[4]), .IN4(n4), .Q(data_o[4]) );
  AO22X1 U10 ( .IN1(data1[3]), .IN2(n5), .IN3(data0[3]), .IN4(n4), .Q(
        data_o[3]) );
  AO22X1 U11 ( .IN1(data1[2]), .IN2(n5), .IN3(data0[2]), .IN4(n4), .Q(
        data_o[2]) );
  AO22X1 U12 ( .IN1(data1[1]), .IN2(n5), .IN3(data0[1]), .IN4(n4), .Q(
        data_o[1]) );
  AO22X1 U13 ( .IN1(data1[15]), .IN2(n5), .IN3(data0[15]), .IN4(n4), .Q(
        data_o[15]) );
  AO22X1 U14 ( .IN1(data1[14]), .IN2(n5), .IN3(data0[14]), .IN4(n4), .Q(
        data_o[14]) );
  AO22X1 U15 ( .IN1(data1[13]), .IN2(n5), .IN3(data0[13]), .IN4(n4), .Q(
        data_o[13]) );
  AO22X1 U16 ( .IN1(data1[12]), .IN2(n5), .IN3(data0[12]), .IN4(n4), .Q(
        data_o[12]) );
  AO22X1 U17 ( .IN1(data1[11]), .IN2(n5), .IN3(data0[11]), .IN4(n4), .Q(
        data_o[11]) );
  AO22X1 U18 ( .IN1(data1[10]), .IN2(n5), .IN3(data0[10]), .IN4(n4), .Q(
        data_o[10]) );
  AO22X1 U19 ( .IN1(data1[0]), .IN2(n5), .IN3(data0[0]), .IN4(n4), .Q(
        data_o[0]) );
  INVX0 U2 ( .INP(select1), .ZN(n1) );
  AND2X1 U3 ( .IN1(select0), .IN2(n1), .Q(n4) );
  NOR2X0 U20 ( .IN1(n1), .IN2(select0), .QN(n5) );
endmodule


module mux3_1_1 ( data0, data1, data2, select0, select1, select2, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  output [15:0] data_o;
  input select0, select1, select2;
  wire   n1, n2, n6, n7, n8;

  AO222X1 U4 ( .IN1(data1[9]), .IN2(n8), .IN3(data0[9]), .IN4(n7), .IN5(
        data2[9]), .IN6(n6), .Q(data_o[9]) );
  AO222X1 U5 ( .IN1(data1[8]), .IN2(n8), .IN3(data0[8]), .IN4(n7), .IN5(
        data2[8]), .IN6(n6), .Q(data_o[8]) );
  AO222X1 U6 ( .IN1(data1[7]), .IN2(n8), .IN3(data0[7]), .IN4(n7), .IN5(
        data2[7]), .IN6(n6), .Q(data_o[7]) );
  AO222X1 U7 ( .IN1(data1[6]), .IN2(n8), .IN3(data0[6]), .IN4(n7), .IN5(
        data2[6]), .IN6(n6), .Q(data_o[6]) );
  AO222X1 U8 ( .IN1(data1[5]), .IN2(n8), .IN3(data0[5]), .IN4(n7), .IN5(
        data2[5]), .IN6(n6), .Q(data_o[5]) );
  AO222X1 U9 ( .IN1(data1[4]), .IN2(n8), .IN3(data0[4]), .IN4(n7), .IN5(
        data2[4]), .IN6(n6), .Q(data_o[4]) );
  AO222X1 U10 ( .IN1(data1[3]), .IN2(n8), .IN3(data0[3]), .IN4(n7), .IN5(
        data2[3]), .IN6(n6), .Q(data_o[3]) );
  AO222X1 U11 ( .IN1(data1[2]), .IN2(n8), .IN3(data0[2]), .IN4(n7), .IN5(
        data2[2]), .IN6(n6), .Q(data_o[2]) );
  AO222X1 U12 ( .IN1(data1[1]), .IN2(n8), .IN3(data0[1]), .IN4(n7), .IN5(
        data2[1]), .IN6(n6), .Q(data_o[1]) );
  AO222X1 U13 ( .IN1(data1[15]), .IN2(n8), .IN3(data0[15]), .IN4(n7), .IN5(
        data2[15]), .IN6(n6), .Q(data_o[15]) );
  AO222X1 U14 ( .IN1(data1[14]), .IN2(n8), .IN3(data0[14]), .IN4(n7), .IN5(
        data2[14]), .IN6(n6), .Q(data_o[14]) );
  AO222X1 U15 ( .IN1(data1[13]), .IN2(n8), .IN3(data0[13]), .IN4(n7), .IN5(
        data2[13]), .IN6(n6), .Q(data_o[13]) );
  AO222X1 U16 ( .IN1(data1[12]), .IN2(n8), .IN3(data0[12]), .IN4(n7), .IN5(
        data2[12]), .IN6(n6), .Q(data_o[12]) );
  AO222X1 U17 ( .IN1(data1[11]), .IN2(n8), .IN3(data0[11]), .IN4(n7), .IN5(
        data2[11]), .IN6(n6), .Q(data_o[11]) );
  AO222X1 U18 ( .IN1(data1[10]), .IN2(n8), .IN3(data0[10]), .IN4(n7), .IN5(
        data2[10]), .IN6(n6), .Q(data_o[10]) );
  AO222X1 U19 ( .IN1(data1[0]), .IN2(n8), .IN3(data0[0]), .IN4(n7), .IN5(
        data2[0]), .IN6(n6), .Q(data_o[0]) );
  INVX0 U2 ( .INP(select0), .ZN(n2) );
  INVX0 U3 ( .INP(select1), .ZN(n1) );
  AND3X1 U20 ( .IN1(n2), .IN2(n1), .IN3(select2), .Q(n6) );
  NOR3X0 U21 ( .IN1(select1), .IN2(select2), .IN3(n2), .QN(n7) );
  NOR3X0 U22 ( .IN1(select0), .IN2(select2), .IN3(n1), .QN(n8) );
endmodule


module mux3_1_0 ( data0, data1, data2, select0, select1, select2, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  output [15:0] data_o;
  input select0, select1, select2;
  wire   n1, n2, n6, n7, n8;

  AO222X1 U4 ( .IN1(data1[9]), .IN2(n8), .IN3(data0[9]), .IN4(n7), .IN5(
        data2[9]), .IN6(n6), .Q(data_o[9]) );
  AO222X1 U5 ( .IN1(data1[8]), .IN2(n8), .IN3(data0[8]), .IN4(n7), .IN5(
        data2[8]), .IN6(n6), .Q(data_o[8]) );
  AO222X1 U6 ( .IN1(data1[7]), .IN2(n8), .IN3(data0[7]), .IN4(n7), .IN5(
        data2[7]), .IN6(n6), .Q(data_o[7]) );
  AO222X1 U7 ( .IN1(data1[6]), .IN2(n8), .IN3(data0[6]), .IN4(n7), .IN5(
        data2[6]), .IN6(n6), .Q(data_o[6]) );
  AO222X1 U8 ( .IN1(data1[5]), .IN2(n8), .IN3(data0[5]), .IN4(n7), .IN5(
        data2[5]), .IN6(n6), .Q(data_o[5]) );
  AO222X1 U9 ( .IN1(data1[4]), .IN2(n8), .IN3(data0[4]), .IN4(n7), .IN5(
        data2[4]), .IN6(n6), .Q(data_o[4]) );
  AO222X1 U10 ( .IN1(data1[3]), .IN2(n8), .IN3(data0[3]), .IN4(n7), .IN5(
        data2[3]), .IN6(n6), .Q(data_o[3]) );
  AO222X1 U11 ( .IN1(data1[2]), .IN2(n8), .IN3(data0[2]), .IN4(n7), .IN5(
        data2[2]), .IN6(n6), .Q(data_o[2]) );
  AO222X1 U12 ( .IN1(data1[1]), .IN2(n8), .IN3(data0[1]), .IN4(n7), .IN5(
        data2[1]), .IN6(n6), .Q(data_o[1]) );
  AO222X1 U13 ( .IN1(data1[15]), .IN2(n8), .IN3(data0[15]), .IN4(n7), .IN5(
        data2[15]), .IN6(n6), .Q(data_o[15]) );
  AO222X1 U14 ( .IN1(data1[14]), .IN2(n8), .IN3(data0[14]), .IN4(n7), .IN5(
        data2[14]), .IN6(n6), .Q(data_o[14]) );
  AO222X1 U15 ( .IN1(data1[13]), .IN2(n8), .IN3(data0[13]), .IN4(n7), .IN5(
        data2[13]), .IN6(n6), .Q(data_o[13]) );
  AO222X1 U16 ( .IN1(data1[12]), .IN2(n8), .IN3(data0[12]), .IN4(n7), .IN5(
        data2[12]), .IN6(n6), .Q(data_o[12]) );
  AO222X1 U17 ( .IN1(data1[11]), .IN2(n8), .IN3(data0[11]), .IN4(n7), .IN5(
        data2[11]), .IN6(n6), .Q(data_o[11]) );
  AO222X1 U18 ( .IN1(data1[10]), .IN2(n8), .IN3(data0[10]), .IN4(n7), .IN5(
        data2[10]), .IN6(n6), .Q(data_o[10]) );
  AO222X1 U19 ( .IN1(data1[0]), .IN2(n8), .IN3(data0[0]), .IN4(n7), .IN5(
        data2[0]), .IN6(n6), .Q(data_o[0]) );
  INVX0 U2 ( .INP(select0), .ZN(n2) );
  INVX0 U3 ( .INP(select1), .ZN(n1) );
  AND3X1 U20 ( .IN1(n2), .IN2(n1), .IN3(select2), .Q(n6) );
  NOR3X0 U21 ( .IN1(select1), .IN2(select2), .IN3(n2), .QN(n7) );
  NOR3X0 U22 ( .IN1(select0), .IN2(select2), .IN3(n1), .QN(n8) );
endmodule



    module node4_NODE_X3_NODE_Y2I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__I_node_2_node_interface__ ( 
        \clk.clk , \reset.reset , \local_node.clk , 
        \local_node.buffer_full_in , \local_node.buffer_full_out , 
        \local_node.receiving_data , \local_node.sending_data , 
        \local_node.data_in , \local_node.data_out , \node_0.clk , 
        \node_0.buffer_full_in , \node_0.buffer_full_out , 
        \node_0.receiving_data , \node_0.sending_data , \node_0.data_in , 
        \node_0.data_out , \node_1.clk , \node_1.buffer_full_in , 
        \node_1.buffer_full_out , \node_1.receiving_data , 
        \node_1.sending_data , \node_1.data_in , \node_1.data_out , 
        \node_2.clk , \node_2.buffer_full_in , \node_2.buffer_full_out , 
        \node_2.receiving_data , \node_2.sending_data , \node_2.data_in , 
        \node_2.data_out  );
  input [15:0] \local_node.data_in ;
  output [15:0] \local_node.data_out ;
  input [15:0] \node_0.data_in ;
  output [15:0] \node_0.data_out ;
  input [15:0] \node_1.data_in ;
  output [15:0] \node_1.data_out ;
  input [15:0] \node_2.data_in ;
  output [15:0] \node_2.data_out ;
  input \clk.clk , \reset.reset , \local_node.buffer_full_in ,
         \local_node.receiving_data , \node_0.buffer_full_in ,
         \node_0.receiving_data , \node_1.buffer_full_in ,
         \node_1.receiving_data , \node_2.buffer_full_in ,
         \node_2.receiving_data ;
  output \local_node.buffer_full_out , \local_node.sending_data ,
         \node_0.buffer_full_out , \node_0.sending_data ,
         \node_1.buffer_full_out , \node_1.sending_data ,
         \node_2.buffer_full_out , \node_2.sending_data ;
  inout \local_node.clk ,  \node_0.clk ,  \node_1.clk ,  \node_2.clk ;
  wire   \buffer_out[3][15] , \buffer_out[3][14] , \buffer_out[3][13] ,
         \buffer_out[3][12] , \buffer_out[3][11] , \buffer_out[3][10] ,
         \buffer_out[3][9] , \buffer_out[3][8] , \buffer_out[3][7] ,
         \buffer_out[3][6] , \buffer_out[3][5] , \buffer_out[3][4] ,
         \buffer_out[3][3] , \buffer_out[3][2] , \buffer_out[3][1] ,
         \buffer_out[3][0] , \buffer_out[2][15] , \buffer_out[2][14] ,
         \buffer_out[2][13] , \buffer_out[2][12] , \buffer_out[2][11] ,
         \buffer_out[2][10] , \buffer_out[2][9] , \buffer_out[2][8] ,
         \buffer_out[2][7] , \buffer_out[2][6] , \buffer_out[2][5] ,
         \buffer_out[2][4] , \buffer_out[2][3] , \buffer_out[2][2] ,
         \buffer_out[2][1] , \buffer_out[2][0] , \buffer_out[1][15] ,
         \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] ,
         \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] ,
         \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] ,
         \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] ,
         \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] ,
         \buffer_out[0][15] , \buffer_out[0][14] , \buffer_out[0][13] ,
         \buffer_out[0][12] , \buffer_out[0][11] , \buffer_out[0][10] ,
         \buffer_out[0][9] , \buffer_out[0][8] , \buffer_out[0][7] ,
         \buffer_out[0][6] , \buffer_out[0][5] , \buffer_out[0][4] ,
         \buffer_out[0][3] , \buffer_out[0][2] , \buffer_out[0][1] ,
         \buffer_out[0][0] , \next_buffer_out[3][15] ,
         \next_buffer_out[3][14] , \next_buffer_out[3][13] ,
         \next_buffer_out[3][12] , \next_buffer_out[3][11] ,
         \next_buffer_out[3][10] , \next_buffer_out[3][9] ,
         \next_buffer_out[3][8] , \next_buffer_out[3][7] ,
         \next_buffer_out[3][6] , \next_buffer_out[3][5] ,
         \next_buffer_out[3][4] , \next_buffer_out[3][3] ,
         \next_buffer_out[3][2] , \next_buffer_out[3][1] ,
         \next_buffer_out[3][0] , \next_buffer_out[2][15] ,
         \next_buffer_out[2][14] , \next_buffer_out[2][13] ,
         \next_buffer_out[2][12] , \next_buffer_out[2][11] ,
         \next_buffer_out[2][10] , \next_buffer_out[2][9] ,
         \next_buffer_out[2][8] , \next_buffer_out[2][7] ,
         \next_buffer_out[2][6] , \next_buffer_out[2][5] ,
         \next_buffer_out[2][4] , \next_buffer_out[2][3] ,
         \next_buffer_out[2][2] , \next_buffer_out[2][1] ,
         \next_buffer_out[2][0] , \next_buffer_out[1][15] ,
         \next_buffer_out[1][14] , \next_buffer_out[1][13] ,
         \next_buffer_out[1][12] , \next_buffer_out[1][11] ,
         \next_buffer_out[1][10] , \next_buffer_out[1][9] ,
         \next_buffer_out[1][8] , \next_buffer_out[1][7] ,
         \next_buffer_out[1][6] , \next_buffer_out[1][5] ,
         \next_buffer_out[1][4] , \next_buffer_out[1][3] ,
         \next_buffer_out[1][2] , \next_buffer_out[1][1] ,
         \next_buffer_out[1][0] , \next_buffer_out[0][15] ,
         \next_buffer_out[0][14] , \next_buffer_out[0][13] ,
         \next_buffer_out[0][12] , \next_buffer_out[0][11] ,
         \next_buffer_out[0][10] , \next_buffer_out[0][9] ,
         \next_buffer_out[0][8] , \next_buffer_out[0][7] ,
         \next_buffer_out[0][6] , \next_buffer_out[0][5] ,
         \next_buffer_out[0][4] , \next_buffer_out[0][3] ,
         \next_buffer_out[0][2] , \next_buffer_out[0][1] ,
         \next_buffer_out[0][0] ;
  wire   [3:0] buffer_full_in;
  wire   [3:0] receiving_data;
  wire   [3:0] pop_v;
  wire   [3:0] data_valid;
  wire   [3:0] next_data_valid;
  wire   [1:0] grant_0;
  wire   [1:0] grant_1;
  wire   [2:0] grant_2;
  wire   [2:0] grant_3;
  tri   \local_node.buffer_full_in ;
  tri   \local_node.buffer_full_out ;
  tri   \local_node.receiving_data ;
  tri   \local_node.sending_data ;
  tri   [15:0] \local_node.data_in ;
  tri   [15:0] \local_node.data_out ;

  converter_out_I_n_node_interface_dut_ c3 ( .\n.buffer_full_in (
        \local_node.buffer_full_in ), .\n.receiving_data (
        \local_node.receiving_data ), .\n.data_in (\local_node.data_in ), 
        .\n.buffer_full_out (\local_node.buffer_full_out ), .\n.sending_data (
        \local_node.sending_data ), .\n.data_out (\local_node.data_out ), 
        .buffer_full_in(1'b0), .receiving_data(1'b0), .data_in({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  fifo_kev_23 \genblk1[0].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[0]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[0]), .data_out({\buffer_out[0][15] , 
        \buffer_out[0][14] , \buffer_out[0][13] , \buffer_out[0][12] , 
        \buffer_out[0][11] , \buffer_out[0][10] , \buffer_out[0][9] , 
        \buffer_out[0][8] , \buffer_out[0][7] , \buffer_out[0][6] , 
        \buffer_out[0][5] , \buffer_out[0][4] , \buffer_out[0][3] , 
        \buffer_out[0][2] , \buffer_out[0][1] , \buffer_out[0][0] }), 
        .next_data_out({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] , 
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .next_data_valid(
        next_data_valid[0]) );
  address_counter_23 \genblk1[0].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] }), 
        .buffer_data_valid(next_data_valid[0]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .buffer_pop(
        pop_v[0]), .receiving_data(1'b0) );
  fifo_kev_22 \genblk1[1].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[1]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[1]), .data_out({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), 
        .next_data_out({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] , 
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .next_data_valid(
        next_data_valid[1]) );
  address_counter_22 \genblk1[1].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] }), 
        .buffer_data_valid(next_data_valid[1]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .buffer_pop(
        pop_v[1]), .receiving_data(1'b0) );
  fifo_kev_21 \genblk1[2].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[2]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[2]), .data_out({\buffer_out[2][15] , 
        \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] , 
        \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] , 
        \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] , 
        \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] , 
        \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] }), 
        .next_data_out({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] , 
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .next_data_valid(
        next_data_valid[2]) );
  address_counter_21 \genblk1[2].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] }), 
        .buffer_data_valid(next_data_valid[2]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .buffer_pop(
        pop_v[2]), .receiving_data(1'b0) );
  fifo_kev_20 \genblk1[3].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[3]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[3]), .data_out({\buffer_out[3][15] , 
        \buffer_out[3][14] , \buffer_out[3][13] , \buffer_out[3][12] , 
        \buffer_out[3][11] , \buffer_out[3][10] , \buffer_out[3][9] , 
        \buffer_out[3][8] , \buffer_out[3][7] , \buffer_out[3][6] , 
        \buffer_out[3][5] , \buffer_out[3][4] , \buffer_out[3][3] , 
        \buffer_out[3][2] , \buffer_out[3][1] , \buffer_out[3][0] }), 
        .next_data_out({\next_buffer_out[3][15] , \next_buffer_out[3][14] , 
        \next_buffer_out[3][13] , \next_buffer_out[3][12] , 
        \next_buffer_out[3][11] , \next_buffer_out[3][10] , 
        \next_buffer_out[3][9] , \next_buffer_out[3][8] , 
        \next_buffer_out[3][7] , \next_buffer_out[3][6] , 
        \next_buffer_out[3][5] , \next_buffer_out[3][4] , 
        \next_buffer_out[3][3] , \next_buffer_out[3][2] , 
        \next_buffer_out[3][1] , \next_buffer_out[3][0] }), .next_data_valid(
        next_data_valid[3]) );
  address_counter_20 \genblk1[3].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[3][15] , \next_buffer_out[3][14] , 
        \next_buffer_out[3][13] , \next_buffer_out[3][12] , 
        \next_buffer_out[3][11] , \next_buffer_out[3][10] , 
        \next_buffer_out[3][9] , \next_buffer_out[3][8] }), 
        .buffer_data_valid(next_data_valid[3]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[3][7] , \next_buffer_out[3][6] , 
        \next_buffer_out[3][5] , \next_buffer_out[3][4] , 
        \next_buffer_out[3][3] , \next_buffer_out[3][2] , 
        \next_buffer_out[3][1] , \next_buffer_out[3][0] }), .buffer_pop(
        pop_v[3]), .receiving_data(1'b0) );
  converter_in_I_n_node_interface_dut__8 \genblk2.c0  ( .\n.buffer_full_in (
        \node_0.buffer_full_in ), .\n.receiving_data (\node_0.receiving_data ), 
        .\n.data_in (\node_0.data_in ), .\n.buffer_full_out (
        \node_0.buffer_full_out ), .\n.sending_data (\node_0.sending_data ), 
        .\n.data_out (\node_0.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_out_I_n_node_interface_dut_ \genblk2.c1  ( .\n.buffer_full_in (
        \node_1.buffer_full_in ), .\n.receiving_data (\node_1.receiving_data ), 
        .\n.data_in (\node_1.data_in ), .\n.buffer_full_out (
        \node_1.buffer_full_out ), .\n.sending_data (\node_1.sending_data ), 
        .\n.data_out (\node_1.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_out_I_n_node_interface_dut_ \genblk2.c2  ( .\n.buffer_full_in (
        \node_2.buffer_full_in ), .\n.receiving_data (\node_2.receiving_data ), 
        .\n.data_in (\node_2.data_in ), .\n.buffer_full_out (
        \node_2.buffer_full_out ), .\n.sending_data (\node_2.sending_data ), 
        .\n.data_out (\node_2.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  controller4_edge_e_0 \genblk2.e  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .packet_addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .local_addr({1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0}), 
        .packet_valid(data_valid), .buffer_full_in({1'b0, 1'b0, 1'b0, 1'b0}), 
        .grant_0(grant_0), .grant_1(grant_1), .grant_2(grant_2), .grant_3(
        grant_3), .pop_v(pop_v) );
  mux2_1_9 \genblk2.mux_n  ( .data0({\buffer_out[1][15] , \buffer_out[1][14] , 
        \buffer_out[1][13] , \buffer_out[1][12] , \buffer_out[1][11] , 
        \buffer_out[1][10] , \buffer_out[1][9] , \buffer_out[1][8] , 
        \buffer_out[1][7] , \buffer_out[1][6] , \buffer_out[1][5] , 
        \buffer_out[1][4] , \buffer_out[1][3] , \buffer_out[1][2] , 
        \buffer_out[1][1] , \buffer_out[1][0] }), .data1({\buffer_out[3][15] , 
        \buffer_out[3][14] , \buffer_out[3][13] , \buffer_out[3][12] , 
        \buffer_out[3][11] , \buffer_out[3][10] , \buffer_out[3][9] , 
        \buffer_out[3][8] , \buffer_out[3][7] , \buffer_out[3][6] , 
        \buffer_out[3][5] , \buffer_out[3][4] , \buffer_out[3][3] , 
        \buffer_out[3][2] , \buffer_out[3][1] , \buffer_out[3][0] }), 
        .select0(grant_0[0]), .select1(grant_0[1]) );
  mux2_1_8 \genblk2.mux_s  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[3][15] , 
        \buffer_out[3][14] , \buffer_out[3][13] , \buffer_out[3][12] , 
        \buffer_out[3][11] , \buffer_out[3][10] , \buffer_out[3][9] , 
        \buffer_out[3][8] , \buffer_out[3][7] , \buffer_out[3][6] , 
        \buffer_out[3][5] , \buffer_out[3][4] , \buffer_out[3][3] , 
        \buffer_out[3][2] , \buffer_out[3][1] , \buffer_out[3][0] }), 
        .select0(grant_1[0]), .select1(grant_1[1]) );
  mux3_1_1 \genblk2.mux_w  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[3][15] , \buffer_out[3][14] , \buffer_out[3][13] , 
        \buffer_out[3][12] , \buffer_out[3][11] , \buffer_out[3][10] , 
        \buffer_out[3][9] , \buffer_out[3][8] , \buffer_out[3][7] , 
        \buffer_out[3][6] , \buffer_out[3][5] , \buffer_out[3][4] , 
        \buffer_out[3][3] , \buffer_out[3][2] , \buffer_out[3][1] , 
        \buffer_out[3][0] }), .select0(grant_2[0]), .select1(grant_2[1]), 
        .select2(grant_2[2]) );
  mux3_1_0 \genblk2.mux_l  ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[2][15] , \buffer_out[2][14] , \buffer_out[2][13] , 
        \buffer_out[2][12] , \buffer_out[2][11] , \buffer_out[2][10] , 
        \buffer_out[2][9] , \buffer_out[2][8] , \buffer_out[2][7] , 
        \buffer_out[2][6] , \buffer_out[2][5] , \buffer_out[2][4] , 
        \buffer_out[2][3] , \buffer_out[2][2] , \buffer_out[2][1] , 
        \buffer_out[2][0] }), .select0(grant_3[0]), .select1(grant_3[1]), 
        .select2(grant_3[2]) );
endmodule


module converter_in_I_n_node_interface_dut__7 ( \n.buffer_full_in , 
        \n.receiving_data , \n.data_in , \n.buffer_full_out , \n.sending_data , 
        \n.data_out , buffer_full_out, sending_data, data_out, buffer_full_in, 
        receiving_data, data_in );
  input [15:0] \n.data_in ;
  output [15:0] \n.data_out ;
  output [15:0] data_out;
  input [15:0] data_in;
  input \n.buffer_full_in , \n.receiving_data , buffer_full_in, receiving_data;
  output \n.buffer_full_out , \n.sending_data , buffer_full_out, sending_data;
  wire   \n.buffer_full_in , \n.receiving_data , buffer_full_in,
         receiving_data;
  assign buffer_full_out = \n.buffer_full_in ;
  assign sending_data = \n.receiving_data ;
  assign data_out[15] = \n.data_in  [15];
  assign data_out[14] = \n.data_in  [14];
  assign data_out[13] = \n.data_in  [13];
  assign data_out[12] = \n.data_in  [12];
  assign data_out[11] = \n.data_in  [11];
  assign data_out[10] = \n.data_in  [10];
  assign data_out[9] = \n.data_in  [9];
  assign data_out[8] = \n.data_in  [8];
  assign data_out[7] = \n.data_in  [7];
  assign data_out[6] = \n.data_in  [6];
  assign data_out[5] = \n.data_in  [5];
  assign data_out[4] = \n.data_in  [4];
  assign data_out[3] = \n.data_in  [3];
  assign data_out[2] = \n.data_in  [2];
  assign data_out[1] = \n.data_in  [1];
  assign data_out[0] = \n.data_in  [0];
  assign \n.buffer_full_out  = buffer_full_in;
  assign \n.sending_data  = receiving_data;
  assign \n.data_out  [15] = data_in[15];
  assign \n.data_out  [14] = data_in[14];
  assign \n.data_out  [13] = data_in[13];
  assign \n.data_out  [12] = data_in[12];
  assign \n.data_out  [11] = data_in[11];
  assign \n.data_out  [10] = data_in[10];
  assign \n.data_out  [9] = data_in[9];
  assign \n.data_out  [8] = data_in[8];
  assign \n.data_out  [7] = data_in[7];
  assign \n.data_out  [6] = data_in[6];
  assign \n.data_out  [5] = data_in[5];
  assign \n.data_out  [4] = data_in[4];
  assign \n.data_out  [3] = data_in[3];
  assign \n.data_out  [2] = data_in[2];
  assign \n.data_out  [1] = data_in[1];
  assign \n.data_out  [0] = data_in[0];

endmodule


module converter_in_I_n_node_interface_dut__6 ( \n.buffer_full_in , 
        \n.receiving_data , \n.data_in , \n.buffer_full_out , \n.sending_data , 
        \n.data_out , buffer_full_out, sending_data, data_out, buffer_full_in, 
        receiving_data, data_in );
  input [15:0] \n.data_in ;
  output [15:0] \n.data_out ;
  output [15:0] data_out;
  input [15:0] data_in;
  input \n.buffer_full_in , \n.receiving_data , buffer_full_in, receiving_data;
  output \n.buffer_full_out , \n.sending_data , buffer_full_out, sending_data;
  wire   \n.buffer_full_in , \n.receiving_data , buffer_full_in,
         receiving_data;
  assign buffer_full_out = \n.buffer_full_in ;
  assign sending_data = \n.receiving_data ;
  assign data_out[15] = \n.data_in  [15];
  assign data_out[14] = \n.data_in  [14];
  assign data_out[13] = \n.data_in  [13];
  assign data_out[12] = \n.data_in  [12];
  assign data_out[11] = \n.data_in  [11];
  assign data_out[10] = \n.data_in  [10];
  assign data_out[9] = \n.data_in  [9];
  assign data_out[8] = \n.data_in  [8];
  assign data_out[7] = \n.data_in  [7];
  assign data_out[6] = \n.data_in  [6];
  assign data_out[5] = \n.data_in  [5];
  assign data_out[4] = \n.data_in  [4];
  assign data_out[3] = \n.data_in  [3];
  assign data_out[2] = \n.data_in  [2];
  assign data_out[1] = \n.data_in  [1];
  assign data_out[0] = \n.data_in  [0];
  assign \n.buffer_full_out  = buffer_full_in;
  assign \n.sending_data  = receiving_data;
  assign \n.data_out  [15] = data_in[15];
  assign \n.data_out  [14] = data_in[14];
  assign \n.data_out  [13] = data_in[13];
  assign \n.data_out  [12] = data_in[12];
  assign \n.data_out  [11] = data_in[11];
  assign \n.data_out  [10] = data_in[10];
  assign \n.data_out  [9] = data_in[9];
  assign \n.data_out  [8] = data_in[8];
  assign \n.data_out  [7] = data_in[7];
  assign \n.data_out  [6] = data_in[6];
  assign \n.data_out  [5] = data_in[5];
  assign \n.data_out  [4] = data_in[4];
  assign \n.data_out  [3] = data_in[3];
  assign \n.data_out  [2] = data_in[2];
  assign \n.data_out  [1] = data_in[1];
  assign \n.data_out  [0] = data_in[0];

endmodule


module fifo_kev_19 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_39 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_19 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_39 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_38 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_19 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_38 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_19_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_19 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_19 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_19 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_19_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_18 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_37 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_18 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_37 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_36 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_18 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_36 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_18_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_18 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_18 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_18 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_18_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_17 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_35 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_17 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_35 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_34 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_17 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_34 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_17_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_17 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_17 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_17 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_17_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_16 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_33 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_16 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_33 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_32 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_16 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_32 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_16_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_16 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_16 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_16 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_16_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_15 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_31 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_15 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_31 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_30 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_15 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_30 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_15_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_15 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_15 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_15 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_15_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module flipflop_BITS2_7 ( clk, data_i, data_o );
  input [1:0] data_i;
  output [1:0] data_o;
  input clk;


  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS2_7 ( clk, enable_i, reset, data_i, data_o );
  input [1:0] data_i;
  input [1:0] data_o;
  input clk, enable_i, reset;
  wire   n10, n11, n1, n5, n7, n8, n9;
  wire   [1:0] write_data;

  AOI22X1 U5 ( .IN1(enable_i), .IN2(data_i[1]), .IN3(n10), .IN4(n1), .QN(n9)
         );
  AOI22X1 U6 ( .IN1(data_i[0]), .IN2(enable_i), .IN3(n11), .IN4(n1), .QN(n8)
         );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n9), .QN(write_data[1]) );
  NOR2X0 U4 ( .IN1(reset), .IN2(n8), .QN(write_data[0]) );
  AND2X1 U7 ( .IN1(data_o[1]), .IN2(n7), .Q(n10) );
  AND2X1 U8 ( .IN1(data_o[0]), .IN2(n5), .Q(n11) );
  flipflop_BITS2_7 FF ( .clk(clk), .data_i(write_data), .data_o({n7, n5}) );
endmodule


module flipflop_BITS1_31 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_31 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_31 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter2_7 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [1:0] request;
  output [1:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   tail_en, n1, n2;
  wire   [1:0] req_i;
  wire   [1:0] req_o;

  AND3X1 U10 ( .IN1(request[1]), .IN2(n1), .IN3(n2), .Q(grant[1]) );
  AND3X1 U11 ( .IN1(request[0]), .IN2(n2), .IN3(request[1]), .Q(tail_en) );
  INVX0 U6 ( .INP(request[0]), .ZN(n1) );
  NOR2X0 U7 ( .IN1(buffer_full_i), .IN2(n1), .QN(grant[0]) );
  INVX0 U8 ( .INP(buffer_full_i), .ZN(n2) );
  OA21X1 U9 ( .IN1(request[1]), .IN2(request[0]), .IN3(n2), .Q(grant_v_o) );
  register_BITS2_7 req_record ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i({1'b1, 1'b0}), .data_o({1'b0, 1'b0}) );
  register_BITS1_31 tail ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i(1'b1), .data_o(1'b0) );
endmodule


module flipflop_BITS2_6 ( clk, data_i, data_o );
  input [1:0] data_i;
  output [1:0] data_o;
  input clk;


  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS2_6 ( clk, enable_i, reset, data_i, data_o );
  input [1:0] data_i;
  input [1:0] data_o;
  input clk, enable_i, reset;
  wire   n10, n11, n1, n5, n7, n8, n9;
  wire   [1:0] write_data;

  AOI22X1 U5 ( .IN1(enable_i), .IN2(data_i[1]), .IN3(n10), .IN4(n1), .QN(n9)
         );
  AOI22X1 U6 ( .IN1(data_i[0]), .IN2(enable_i), .IN3(n11), .IN4(n1), .QN(n8)
         );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n9), .QN(write_data[1]) );
  NOR2X0 U4 ( .IN1(reset), .IN2(n8), .QN(write_data[0]) );
  AND2X1 U7 ( .IN1(data_o[1]), .IN2(n7), .Q(n10) );
  AND2X1 U8 ( .IN1(data_o[0]), .IN2(n5), .Q(n11) );
  flipflop_BITS2_6 FF ( .clk(clk), .data_i(write_data), .data_o({n7, n5}) );
endmodule


module flipflop_BITS1_30 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_30 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_30 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter2_6 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [1:0] request;
  output [1:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   tail_en, n1, n2;
  wire   [1:0] req_i;
  wire   [1:0] req_o;

  AND3X1 U10 ( .IN1(request[1]), .IN2(n1), .IN3(n2), .Q(grant[1]) );
  AND3X1 U11 ( .IN1(request[0]), .IN2(n2), .IN3(request[1]), .Q(tail_en) );
  INVX0 U6 ( .INP(request[0]), .ZN(n1) );
  NOR2X0 U7 ( .IN1(buffer_full_i), .IN2(n1), .QN(grant[0]) );
  INVX0 U8 ( .INP(buffer_full_i), .ZN(n2) );
  OA21X1 U9 ( .IN1(request[1]), .IN2(request[0]), .IN3(n2), .Q(grant_v_o) );
  register_BITS2_6 req_record ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i({1'b1, 1'b0}), .data_o({1'b0, 1'b0}) );
  register_BITS1_30 tail ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i(1'b1), .data_o(1'b0) );
endmodule


module flipflop_BITS4_35 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_35 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_35 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS4_34 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_34 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_34 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS4_33 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_33 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_33 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS1_29 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_29 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_29 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_28 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_28 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_28 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter4_11 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [3:0] request;
  output [3:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[2][3] , \req_i[2][2] , \req_i[2][1] , \req_i[2][0] ,
         \req_i[1][3] , \req_i[1][2] , \req_i[1][1] , \req_i[1][0] ,
         \req_i[0][3] , \req_i[0][2] , \req_i[0][1] , tail_en, N71, N265, N266,
         N267, N268, N276, N282, N291, N300, N301, N302, N303, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n1, n2, n3, n4, n6,
         n7;
  wire   [2:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N265 = request[0];
  assign N266 = request[1];
  assign N267 = request[2];
  assign N268 = request[3];

  LATCHX1 shift_reg ( .CLK(1'b0), .D(1'b0), .Q(N71) );
  LATCHX1 \grant_reg[3]  ( .CLK(1'b1), .D(N303), .Q(grant[3]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N302), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N301), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N300), .Q(grant[0]) );
  LNANDX1 \req_i_reg[2][3]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][3] ) );
  LNANDX1 \req_i_reg[2][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][2] ) );
  LNANDX1 \req_i_reg[2][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][1] ) );
  LNANDX1 \req_i_reg[2][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][0] ) );
  LNANDX1 \req_i_reg[1][3]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][3] ) );
  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][3]  ( .CLK(tail_en), .D(N282), .Q(\req_i[0][3] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(n1), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(n4), .Q(\req_i[0][1] ) );
  LATCHX1 \tail_i_reg[0]  ( .CLK(tail_en), .D(N276), .Q(tail_i[0]) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N291), .D(tail_en), .Q(req_en[0]) );
  AND3X1 U35 ( .IN1(grant_v_o), .IN2(n72), .IN3(N267), .Q(N302) );
  NAND4X0 U37 ( .IN1(n74), .IN2(grant_v_o), .IN3(n75), .IN4(n71), .QN(N291) );
  AO21X1 U38 ( .IN1(n77), .IN2(n72), .IN3(buffer_full_i), .Q(n70) );
  NOR3X0 U39 ( .IN1(n4), .IN2(N282), .IN3(n1), .QN(n74) );
  NAND4X0 U41 ( .IN1(n80), .IN2(n78), .IN3(n82), .IN4(n81), .QN(N276) );
  AOI22X1 U42 ( .IN1(n2), .IN2(n76), .IN3(n76), .IN4(N265), .QN(n78) );
  AND2X1 U43 ( .IN1(N268), .IN2(n6), .Q(n76) );
  OA22X1 U44 ( .IN1(n6), .IN2(n73), .IN3(n6), .IN4(n3), .Q(n80) );
  INVX0 U15 ( .INP(N267), .ZN(n6) );
  INVX0 U16 ( .INP(n73), .ZN(n2) );
  NAND2X1 U17 ( .IN1(N266), .IN2(N265), .QN(n81) );
  NAND2X1 U18 ( .IN1(N267), .IN2(N268), .QN(n79) );
  INVX0 U19 ( .INP(N265), .ZN(n3) );
  NAND2X1 U20 ( .IN1(N266), .IN2(n3), .QN(n73) );
  NOR2X0 U21 ( .IN1(N266), .IN2(N265), .QN(n72) );
  INVX0 U22 ( .INP(n70), .ZN(grant_v_o) );
  NOR2X0 U23 ( .IN1(N268), .IN2(N267), .QN(n77) );
  NAND2X1 U24 ( .IN1(n76), .IN2(n72), .QN(n71) );
  NOR2X0 U25 ( .IN1(N265), .IN2(n2), .QN(n75) );
  NAND2X1 U26 ( .IN1(N71), .IN2(n7), .QN(n82) );
  INVX0 U27 ( .INP(n79), .ZN(n7) );
  INVX0 U28 ( .INP(n81), .ZN(n4) );
  INVX0 U29 ( .INP(n80), .ZN(n1) );
  NAND2X1 U30 ( .IN1(n78), .IN2(n79), .QN(N282) );
  NOR2X0 U31 ( .IN1(n70), .IN2(n74), .QN(tail_en) );
  NOR2X0 U32 ( .IN1(n3), .IN2(n70), .QN(N300) );
  NOR2X0 U33 ( .IN1(n73), .IN2(n70), .QN(N301) );
  NOR2X0 U34 ( .IN1(n70), .IN2(n71), .QN(N303) );
  register_BITS4_35 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][3] , \req_i[0][2] , \req_i[0][1] , 
        1'b0}), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS4_34 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][3] , \req_i[1][2] , \req_i[1][1] , 
        \req_i[1][0] }), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS4_33 \genblk1[2].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[2][3] , \req_i[2][2] , \req_i[2][1] , 
        \req_i[2][0] }), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS1_29 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(tail_i[0]), .data_o(1'b0) );
  register_BITS1_28 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module flipflop_BITS4_32 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_32 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_32 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS4_31 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_31 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_31 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS4_30 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_30 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_30 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS1_27 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_27 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_27 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_26 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_26 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_26 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter4_10 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [3:0] request;
  output [3:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[2][3] , \req_i[2][2] , \req_i[2][1] , \req_i[2][0] ,
         \req_i[1][3] , \req_i[1][2] , \req_i[1][1] , \req_i[1][0] ,
         \req_i[0][3] , \req_i[0][2] , \req_i[0][1] , tail_en, N71, N265, N266,
         N267, N268, N276, N282, N291, N300, N301, N302, N303, n1, n2, n3, n4,
         n6, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21;
  wire   [2:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N265 = request[0];
  assign N266 = request[1];
  assign N267 = request[2];
  assign N268 = request[3];

  LATCHX1 shift_reg ( .CLK(1'b0), .D(1'b0), .Q(N71) );
  LATCHX1 \grant_reg[3]  ( .CLK(1'b1), .D(N303), .Q(grant[3]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N302), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N301), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N300), .Q(grant[0]) );
  LNANDX1 \req_i_reg[2][3]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][3] ) );
  LNANDX1 \req_i_reg[2][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][2] ) );
  LNANDX1 \req_i_reg[2][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][1] ) );
  LNANDX1 \req_i_reg[2][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][0] ) );
  LNANDX1 \req_i_reg[1][3]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][3] ) );
  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][3]  ( .CLK(tail_en), .D(N282), .Q(\req_i[0][3] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(n1), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(n4), .Q(\req_i[0][1] ) );
  LATCHX1 \tail_i_reg[0]  ( .CLK(tail_en), .D(N276), .Q(tail_i[0]) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N291), .D(tail_en), .Q(req_en[0]) );
  AND3X1 U35 ( .IN1(grant_v_o), .IN2(n19), .IN3(N267), .Q(N302) );
  NAND4X0 U37 ( .IN1(n17), .IN2(grant_v_o), .IN3(n16), .IN4(n20), .QN(N291) );
  AO21X1 U38 ( .IN1(n14), .IN2(n19), .IN3(buffer_full_i), .Q(n21) );
  NOR3X0 U39 ( .IN1(n4), .IN2(N282), .IN3(n1), .QN(n17) );
  NAND4X0 U41 ( .IN1(n11), .IN2(n13), .IN3(n9), .IN4(n10), .QN(N276) );
  AOI22X1 U42 ( .IN1(n2), .IN2(n15), .IN3(n15), .IN4(N265), .QN(n13) );
  AND2X1 U43 ( .IN1(N268), .IN2(n6), .Q(n15) );
  OA22X1 U44 ( .IN1(n6), .IN2(n18), .IN3(n6), .IN4(n3), .Q(n11) );
  INVX0 U15 ( .INP(N267), .ZN(n6) );
  INVX0 U16 ( .INP(n18), .ZN(n2) );
  NAND2X1 U17 ( .IN1(N266), .IN2(N265), .QN(n10) );
  NAND2X1 U18 ( .IN1(N267), .IN2(N268), .QN(n12) );
  INVX0 U19 ( .INP(N265), .ZN(n3) );
  NAND2X1 U20 ( .IN1(N266), .IN2(n3), .QN(n18) );
  NOR2X0 U21 ( .IN1(N266), .IN2(N265), .QN(n19) );
  INVX0 U22 ( .INP(n21), .ZN(grant_v_o) );
  NOR2X0 U23 ( .IN1(N268), .IN2(N267), .QN(n14) );
  NAND2X1 U24 ( .IN1(n15), .IN2(n19), .QN(n20) );
  NOR2X0 U25 ( .IN1(N265), .IN2(n2), .QN(n16) );
  NAND2X1 U26 ( .IN1(N71), .IN2(n7), .QN(n9) );
  INVX0 U27 ( .INP(n12), .ZN(n7) );
  INVX0 U28 ( .INP(n10), .ZN(n4) );
  INVX0 U29 ( .INP(n11), .ZN(n1) );
  NAND2X1 U30 ( .IN1(n13), .IN2(n12), .QN(N282) );
  NOR2X0 U31 ( .IN1(n21), .IN2(n17), .QN(tail_en) );
  NOR2X0 U32 ( .IN1(n3), .IN2(n21), .QN(N300) );
  NOR2X0 U33 ( .IN1(n18), .IN2(n21), .QN(N301) );
  NOR2X0 U34 ( .IN1(n21), .IN2(n20), .QN(N303) );
  register_BITS4_32 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][3] , \req_i[0][2] , \req_i[0][1] , 
        1'b0}), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS4_31 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][3] , \req_i[1][2] , \req_i[1][1] , 
        \req_i[1][0] }), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS4_30 \genblk1[2].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[2][3] , \req_i[2][2] , \req_i[2][1] , 
        \req_i[2][0] }), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS1_27 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(tail_i[0]), .data_o(1'b0) );
  register_BITS1_26 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module flipflop_BITS4_29 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_29 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_29 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS4_28 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_28 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_28 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS4_27 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_27 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_27 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS1_25 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_25 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_25 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_24 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_24 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_24 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter4_9 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [3:0] request;
  output [3:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[2][3] , \req_i[2][2] , \req_i[2][1] , \req_i[2][0] ,
         \req_i[1][3] , \req_i[1][2] , \req_i[1][1] , \req_i[1][0] ,
         \req_i[0][3] , \req_i[0][2] , \req_i[0][1] , tail_en, N71, N265, N266,
         N267, N268, N276, N282, N291, N300, N301, N302, N303, n1, n2, n3, n4,
         n6, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21;
  wire   [2:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N265 = request[0];
  assign N266 = request[1];
  assign N267 = request[2];
  assign N268 = request[3];

  LATCHX1 shift_reg ( .CLK(1'b0), .D(1'b0), .Q(N71) );
  LATCHX1 \grant_reg[3]  ( .CLK(1'b1), .D(N303), .Q(grant[3]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N302), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N301), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N300), .Q(grant[0]) );
  LNANDX1 \req_i_reg[2][3]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][3] ) );
  LNANDX1 \req_i_reg[2][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][2] ) );
  LNANDX1 \req_i_reg[2][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][1] ) );
  LNANDX1 \req_i_reg[2][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][0] ) );
  LNANDX1 \req_i_reg[1][3]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][3] ) );
  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][3]  ( .CLK(tail_en), .D(N282), .Q(\req_i[0][3] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(n1), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(n4), .Q(\req_i[0][1] ) );
  LATCHX1 \tail_i_reg[0]  ( .CLK(tail_en), .D(N276), .Q(tail_i[0]) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N291), .D(tail_en), .Q(req_en[0]) );
  AND3X1 U35 ( .IN1(grant_v_o), .IN2(n19), .IN3(N267), .Q(N302) );
  NAND4X0 U37 ( .IN1(n17), .IN2(grant_v_o), .IN3(n16), .IN4(n20), .QN(N291) );
  AO21X1 U38 ( .IN1(n14), .IN2(n19), .IN3(buffer_full_i), .Q(n21) );
  NOR3X0 U39 ( .IN1(n4), .IN2(N282), .IN3(n1), .QN(n17) );
  NAND4X0 U41 ( .IN1(n11), .IN2(n13), .IN3(n9), .IN4(n10), .QN(N276) );
  AOI22X1 U42 ( .IN1(n2), .IN2(n15), .IN3(n15), .IN4(N265), .QN(n13) );
  AND2X1 U43 ( .IN1(N268), .IN2(n6), .Q(n15) );
  OA22X1 U44 ( .IN1(n6), .IN2(n18), .IN3(n6), .IN4(n3), .Q(n11) );
  INVX0 U15 ( .INP(N267), .ZN(n6) );
  INVX0 U16 ( .INP(n18), .ZN(n2) );
  NAND2X1 U17 ( .IN1(N266), .IN2(N265), .QN(n10) );
  NAND2X1 U18 ( .IN1(N267), .IN2(N268), .QN(n12) );
  INVX0 U19 ( .INP(N265), .ZN(n3) );
  NAND2X1 U20 ( .IN1(N266), .IN2(n3), .QN(n18) );
  NOR2X0 U21 ( .IN1(N266), .IN2(N265), .QN(n19) );
  INVX0 U22 ( .INP(n21), .ZN(grant_v_o) );
  NOR2X0 U23 ( .IN1(N268), .IN2(N267), .QN(n14) );
  NAND2X1 U24 ( .IN1(n15), .IN2(n19), .QN(n20) );
  NOR2X0 U25 ( .IN1(N265), .IN2(n2), .QN(n16) );
  NAND2X1 U26 ( .IN1(N71), .IN2(n7), .QN(n9) );
  INVX0 U27 ( .INP(n12), .ZN(n7) );
  INVX0 U28 ( .INP(n10), .ZN(n4) );
  INVX0 U29 ( .INP(n11), .ZN(n1) );
  NAND2X1 U30 ( .IN1(n13), .IN2(n12), .QN(N282) );
  NOR2X0 U31 ( .IN1(n21), .IN2(n17), .QN(tail_en) );
  NOR2X0 U32 ( .IN1(n3), .IN2(n21), .QN(N300) );
  NOR2X0 U33 ( .IN1(n18), .IN2(n21), .QN(N301) );
  NOR2X0 U34 ( .IN1(n21), .IN2(n20), .QN(N303) );
  register_BITS4_29 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][3] , \req_i[0][2] , \req_i[0][1] , 
        1'b0}), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS4_28 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][3] , \req_i[1][2] , \req_i[1][1] , 
        \req_i[1][0] }), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS4_27 \genblk1[2].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[2][3] , \req_i[2][2] , \req_i[2][1] , 
        \req_i[2][0] }), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS1_25 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(tail_i[0]), .data_o(1'b0) );
  register_BITS1_24 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module dccl_19 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_18 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_17 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_16 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_15 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module controller5_3 ( clk, rst, .packet_addr({\packet_addr[4][7] , 
        \packet_addr[4][6] , \packet_addr[4][5] , \packet_addr[4][4] , 
        \packet_addr[4][3] , \packet_addr[4][2] , \packet_addr[4][1] , 
        \packet_addr[4][0] , \packet_addr[3][7] , \packet_addr[3][6] , 
        \packet_addr[3][5] , \packet_addr[3][4] , \packet_addr[3][3] , 
        \packet_addr[3][2] , \packet_addr[3][1] , \packet_addr[3][0] , 
        \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] , 
        \packet_addr[2][4] , \packet_addr[2][3] , \packet_addr[2][2] , 
        \packet_addr[2][1] , \packet_addr[2][0] , \packet_addr[1][7] , 
        \packet_addr[1][6] , \packet_addr[1][5] , \packet_addr[1][4] , 
        \packet_addr[1][3] , \packet_addr[1][2] , \packet_addr[1][1] , 
        \packet_addr[1][0] , \packet_addr[0][7] , \packet_addr[0][6] , 
        \packet_addr[0][5] , \packet_addr[0][4] , \packet_addr[0][3] , 
        \packet_addr[0][2] , \packet_addr[0][1] , \packet_addr[0][0] }), 
        local_addr, packet_valid, buffer_full_in, grant_0, grant_1, grant_2, 
        grant_3, grant_4, grant_v, pop_v );
  input [7:0] local_addr;
  input [4:0] packet_valid;
  input [4:0] buffer_full_in;
  output [1:0] grant_0;
  output [1:0] grant_1;
  output [3:0] grant_2;
  output [3:0] grant_3;
  output [3:0] grant_4;
  output [4:0] grant_v;
  output [4:0] pop_v;
  input clk, rst, \packet_addr[4][7] , \packet_addr[4][6] ,
         \packet_addr[4][5] , \packet_addr[4][4] , \packet_addr[4][3] ,
         \packet_addr[4][2] , \packet_addr[4][1] , \packet_addr[4][0] ,
         \packet_addr[3][7] , \packet_addr[3][6] , \packet_addr[3][5] ,
         \packet_addr[3][4] , \packet_addr[3][3] , \packet_addr[3][2] ,
         \packet_addr[3][1] , \packet_addr[3][0] , \packet_addr[2][7] ,
         \packet_addr[2][6] , \packet_addr[2][5] , \packet_addr[2][4] ,
         \packet_addr[2][3] , \packet_addr[2][2] , \packet_addr[2][1] ,
         \packet_addr[2][0] , \packet_addr[1][7] , \packet_addr[1][6] ,
         \packet_addr[1][5] , \packet_addr[1][4] , \packet_addr[1][3] ,
         \packet_addr[1][2] , \packet_addr[1][1] , \packet_addr[1][0] ,
         \packet_addr[0][7] , \packet_addr[0][6] , \packet_addr[0][5] ,
         \packet_addr[0][4] , \packet_addr[0][3] , \packet_addr[0][2] ,
         \packet_addr[0][1] , \packet_addr[0][0] ;
  wire   \request[4][3] , \request[4][2] , \request[4][1] , \request[4][0] ,
         \request[3][3] , \request[3][2] , \request[3][1] , \request[3][0] ,
         \request[2][3] , \request[2][2] , \request[2][1] , \request[2][0] ,
         \request[1][1] , \request[1][0] , \request[0][1] , \request[0][0] ;

  OR4X1 U1 ( .IN1(grant_1[1]), .IN2(grant_0[1]), .IN3(grant_3[3]), .IN4(
        grant_2[3]), .Q(pop_v[4]) );
  OR2X1 U2 ( .IN1(grant_2[2]), .IN2(grant_4[3]), .Q(pop_v[3]) );
  OR2X1 U3 ( .IN1(grant_3[2]), .IN2(grant_4[2]), .Q(pop_v[2]) );
  OR4X1 U4 ( .IN1(grant_2[1]), .IN2(grant_0[0]), .IN3(grant_4[1]), .IN4(
        grant_3[1]), .Q(pop_v[1]) );
  OR4X1 U5 ( .IN1(grant_2[0]), .IN2(grant_1[0]), .IN3(grant_4[0]), .IN4(
        grant_3[0]), .Q(pop_v[0]) );
  arbiter2_7 arbiter_n ( .clk(clk), .rst(rst), .request({\request[0][1] , 
        \request[0][0] }), .buffer_full_i(buffer_full_in[0]), .grant(grant_0), 
        .grant_v_o(grant_v[0]) );
  arbiter2_6 arbiter_s ( .clk(clk), .rst(rst), .request({\request[1][1] , 
        \request[1][0] }), .buffer_full_i(buffer_full_in[1]), .grant(grant_1), 
        .grant_v_o(grant_v[1]) );
  arbiter4_11 arbiter_e ( .clk(clk), .rst(rst), .request({\request[2][3] , 
        \request[2][2] , \request[2][1] , \request[2][0] }), .buffer_full_i(
        buffer_full_in[2]), .grant(grant_2), .grant_v_o(grant_v[2]) );
  arbiter4_10 arbiter_w ( .clk(clk), .rst(rst), .request({\request[3][3] , 
        \request[3][2] , \request[3][1] , \request[3][0] }), .buffer_full_i(
        buffer_full_in[3]), .grant(grant_3), .grant_v_o(grant_v[3]) );
  arbiter4_9 arbiter_l ( .clk(clk), .rst(rst), .request({\request[4][3] , 
        \request[4][2] , \request[4][1] , \request[4][0] }), .buffer_full_i(
        buffer_full_in[4]), .grant(grant_4), .grant_v_o(grant_v[4]) );
  dccl_19 dccl_n ( .packet_addr_y_i({\packet_addr[0][3] , \packet_addr[0][2] , 
        \packet_addr[0][1] , \packet_addr[0][0] }), .packet_addr_x_i({
        \packet_addr[0][7] , \packet_addr[0][6] , \packet_addr[0][5] , 
        \packet_addr[0][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[0]), 
        .east_req(\request[2][0] ), .south_req(\request[1][0] ), .west_req(
        \request[3][0] ), .local_req(\request[4][0] ) );
  dccl_18 dccl_s ( .packet_addr_y_i({\packet_addr[1][3] , \packet_addr[1][2] , 
        \packet_addr[1][1] , \packet_addr[1][0] }), .packet_addr_x_i({
        \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] , 
        \packet_addr[1][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[1]), 
        .north_req(\request[0][0] ), .east_req(\request[2][1] ), .west_req(
        \request[3][1] ), .local_req(\request[4][1] ) );
  dccl_17 dccl_e ( .packet_addr_y_i({\packet_addr[2][3] , \packet_addr[2][2] , 
        \packet_addr[2][1] , \packet_addr[2][0] }), .packet_addr_x_i({
        \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] , 
        \packet_addr[2][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[2]), 
        .west_req(\request[3][2] ), .local_req(\request[4][2] ) );
  dccl_16 dccl_w ( .packet_addr_y_i({\packet_addr[3][3] , \packet_addr[3][2] , 
        \packet_addr[3][1] , \packet_addr[3][0] }), .packet_addr_x_i({
        \packet_addr[3][7] , \packet_addr[3][6] , \packet_addr[3][5] , 
        \packet_addr[3][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[3]), 
        .east_req(\request[2][2] ), .local_req(\request[4][3] ) );
  dccl_15 dccl_l ( .packet_addr_y_i({\packet_addr[4][3] , \packet_addr[4][2] , 
        \packet_addr[4][1] , \packet_addr[4][0] }), .packet_addr_x_i({
        \packet_addr[4][7] , \packet_addr[4][6] , \packet_addr[4][5] , 
        \packet_addr[4][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[4]), 
        .north_req(\request[0][1] ), .east_req(\request[2][3] ), .south_req(
        \request[1][1] ), .west_req(\request[3][3] ) );
endmodule


module mux2_1_7 ( data0, data1, select0, select1, data_o );
  input [15:0] data0;
  input [15:0] data1;
  output [15:0] data_o;
  input select0, select1;
  wire   n1, n4, n5;

  AO22X1 U4 ( .IN1(data1[9]), .IN2(n5), .IN3(data0[9]), .IN4(n4), .Q(data_o[9]) );
  AO22X1 U5 ( .IN1(data1[8]), .IN2(n5), .IN3(data0[8]), .IN4(n4), .Q(data_o[8]) );
  AO22X1 U6 ( .IN1(data1[7]), .IN2(n5), .IN3(data0[7]), .IN4(n4), .Q(data_o[7]) );
  AO22X1 U7 ( .IN1(data1[6]), .IN2(n5), .IN3(data0[6]), .IN4(n4), .Q(data_o[6]) );
  AO22X1 U8 ( .IN1(data1[5]), .IN2(n5), .IN3(data0[5]), .IN4(n4), .Q(data_o[5]) );
  AO22X1 U9 ( .IN1(data1[4]), .IN2(n5), .IN3(data0[4]), .IN4(n4), .Q(data_o[4]) );
  AO22X1 U10 ( .IN1(data1[3]), .IN2(n5), .IN3(data0[3]), .IN4(n4), .Q(
        data_o[3]) );
  AO22X1 U11 ( .IN1(data1[2]), .IN2(n5), .IN3(data0[2]), .IN4(n4), .Q(
        data_o[2]) );
  AO22X1 U12 ( .IN1(data1[1]), .IN2(n5), .IN3(data0[1]), .IN4(n4), .Q(
        data_o[1]) );
  AO22X1 U13 ( .IN1(data1[15]), .IN2(n5), .IN3(data0[15]), .IN4(n4), .Q(
        data_o[15]) );
  AO22X1 U14 ( .IN1(data1[14]), .IN2(n5), .IN3(data0[14]), .IN4(n4), .Q(
        data_o[14]) );
  AO22X1 U15 ( .IN1(data1[13]), .IN2(n5), .IN3(data0[13]), .IN4(n4), .Q(
        data_o[13]) );
  AO22X1 U16 ( .IN1(data1[12]), .IN2(n5), .IN3(data0[12]), .IN4(n4), .Q(
        data_o[12]) );
  AO22X1 U17 ( .IN1(data1[11]), .IN2(n5), .IN3(data0[11]), .IN4(n4), .Q(
        data_o[11]) );
  AO22X1 U18 ( .IN1(data1[10]), .IN2(n5), .IN3(data0[10]), .IN4(n4), .Q(
        data_o[10]) );
  AO22X1 U19 ( .IN1(data1[0]), .IN2(n5), .IN3(data0[0]), .IN4(n4), .Q(
        data_o[0]) );
  INVX0 U2 ( .INP(select1), .ZN(n1) );
  AND2X1 U3 ( .IN1(select0), .IN2(n1), .Q(n4) );
  NOR2X0 U20 ( .IN1(n1), .IN2(select0), .QN(n5) );
endmodule


module mux2_1_6 ( data0, data1, select0, select1, data_o );
  input [15:0] data0;
  input [15:0] data1;
  output [15:0] data_o;
  input select0, select1;
  wire   n1, n4, n5;

  AO22X1 U4 ( .IN1(data1[9]), .IN2(n5), .IN3(data0[9]), .IN4(n4), .Q(data_o[9]) );
  AO22X1 U5 ( .IN1(data1[8]), .IN2(n5), .IN3(data0[8]), .IN4(n4), .Q(data_o[8]) );
  AO22X1 U6 ( .IN1(data1[7]), .IN2(n5), .IN3(data0[7]), .IN4(n4), .Q(data_o[7]) );
  AO22X1 U7 ( .IN1(data1[6]), .IN2(n5), .IN3(data0[6]), .IN4(n4), .Q(data_o[6]) );
  AO22X1 U8 ( .IN1(data1[5]), .IN2(n5), .IN3(data0[5]), .IN4(n4), .Q(data_o[5]) );
  AO22X1 U9 ( .IN1(data1[4]), .IN2(n5), .IN3(data0[4]), .IN4(n4), .Q(data_o[4]) );
  AO22X1 U10 ( .IN1(data1[3]), .IN2(n5), .IN3(data0[3]), .IN4(n4), .Q(
        data_o[3]) );
  AO22X1 U11 ( .IN1(data1[2]), .IN2(n5), .IN3(data0[2]), .IN4(n4), .Q(
        data_o[2]) );
  AO22X1 U12 ( .IN1(data1[1]), .IN2(n5), .IN3(data0[1]), .IN4(n4), .Q(
        data_o[1]) );
  AO22X1 U13 ( .IN1(data1[15]), .IN2(n5), .IN3(data0[15]), .IN4(n4), .Q(
        data_o[15]) );
  AO22X1 U14 ( .IN1(data1[14]), .IN2(n5), .IN3(data0[14]), .IN4(n4), .Q(
        data_o[14]) );
  AO22X1 U15 ( .IN1(data1[13]), .IN2(n5), .IN3(data0[13]), .IN4(n4), .Q(
        data_o[13]) );
  AO22X1 U16 ( .IN1(data1[12]), .IN2(n5), .IN3(data0[12]), .IN4(n4), .Q(
        data_o[12]) );
  AO22X1 U17 ( .IN1(data1[11]), .IN2(n5), .IN3(data0[11]), .IN4(n4), .Q(
        data_o[11]) );
  AO22X1 U18 ( .IN1(data1[10]), .IN2(n5), .IN3(data0[10]), .IN4(n4), .Q(
        data_o[10]) );
  AO22X1 U19 ( .IN1(data1[0]), .IN2(n5), .IN3(data0[0]), .IN4(n4), .Q(
        data_o[0]) );
  INVX0 U2 ( .INP(select1), .ZN(n1) );
  AND2X1 U3 ( .IN1(select0), .IN2(n1), .Q(n4) );
  NOR2X0 U20 ( .IN1(n1), .IN2(select0), .QN(n5) );
endmodule


module mux4_1_11 ( data0, data1, data2, data3, select0, select1, select2, 
        select3, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  input [15:0] data3;
  output [15:0] data_o;
  input select0, select1, select2, select3;
  wire   n1, n2, n3, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43;

  AO221X1 U5 ( .IN1(data1[9]), .IN2(n43), .IN3(data0[9]), .IN4(n42), .IN5(n41), 
        .Q(data_o[9]) );
  AO22X1 U6 ( .IN1(data2[9]), .IN2(n40), .IN3(data3[9]), .IN4(n39), .Q(n41) );
  AO221X1 U7 ( .IN1(data1[8]), .IN2(n43), .IN3(data0[8]), .IN4(n42), .IN5(n38), 
        .Q(data_o[8]) );
  AO22X1 U8 ( .IN1(data2[8]), .IN2(n40), .IN3(data3[8]), .IN4(n39), .Q(n38) );
  AO221X1 U9 ( .IN1(data1[7]), .IN2(n43), .IN3(data0[7]), .IN4(n42), .IN5(n37), 
        .Q(data_o[7]) );
  AO22X1 U10 ( .IN1(data2[7]), .IN2(n40), .IN3(data3[7]), .IN4(n39), .Q(n37)
         );
  AO221X1 U11 ( .IN1(data1[6]), .IN2(n43), .IN3(data0[6]), .IN4(n42), .IN5(n36), .Q(data_o[6]) );
  AO22X1 U12 ( .IN1(data2[6]), .IN2(n40), .IN3(data3[6]), .IN4(n39), .Q(n36)
         );
  AO221X1 U13 ( .IN1(data1[5]), .IN2(n43), .IN3(data0[5]), .IN4(n42), .IN5(n35), .Q(data_o[5]) );
  AO22X1 U14 ( .IN1(data2[5]), .IN2(n40), .IN3(data3[5]), .IN4(n39), .Q(n35)
         );
  AO221X1 U15 ( .IN1(data1[4]), .IN2(n43), .IN3(data0[4]), .IN4(n42), .IN5(n34), .Q(data_o[4]) );
  AO22X1 U16 ( .IN1(data2[4]), .IN2(n40), .IN3(data3[4]), .IN4(n39), .Q(n34)
         );
  AO221X1 U17 ( .IN1(data1[3]), .IN2(n43), .IN3(data0[3]), .IN4(n42), .IN5(n33), .Q(data_o[3]) );
  AO22X1 U18 ( .IN1(data2[3]), .IN2(n40), .IN3(data3[3]), .IN4(n39), .Q(n33)
         );
  AO221X1 U19 ( .IN1(data1[2]), .IN2(n43), .IN3(data0[2]), .IN4(n42), .IN5(n32), .Q(data_o[2]) );
  AO22X1 U20 ( .IN1(data2[2]), .IN2(n40), .IN3(data3[2]), .IN4(n39), .Q(n32)
         );
  AO221X1 U21 ( .IN1(data1[1]), .IN2(n43), .IN3(data0[1]), .IN4(n42), .IN5(n31), .Q(data_o[1]) );
  AO22X1 U22 ( .IN1(data2[1]), .IN2(n40), .IN3(data3[1]), .IN4(n39), .Q(n31)
         );
  AO221X1 U23 ( .IN1(data1[15]), .IN2(n43), .IN3(data0[15]), .IN4(n42), .IN5(
        n30), .Q(data_o[15]) );
  AO22X1 U24 ( .IN1(data2[15]), .IN2(n40), .IN3(data3[15]), .IN4(n39), .Q(n30)
         );
  AO221X1 U25 ( .IN1(data1[14]), .IN2(n43), .IN3(data0[14]), .IN4(n42), .IN5(
        n29), .Q(data_o[14]) );
  AO22X1 U26 ( .IN1(data2[14]), .IN2(n40), .IN3(data3[14]), .IN4(n39), .Q(n29)
         );
  AO221X1 U27 ( .IN1(data1[13]), .IN2(n43), .IN3(data0[13]), .IN4(n42), .IN5(
        n28), .Q(data_o[13]) );
  AO22X1 U28 ( .IN1(data2[13]), .IN2(n40), .IN3(data3[13]), .IN4(n39), .Q(n28)
         );
  AO221X1 U29 ( .IN1(data1[12]), .IN2(n43), .IN3(data0[12]), .IN4(n42), .IN5(
        n27), .Q(data_o[12]) );
  AO22X1 U30 ( .IN1(data2[12]), .IN2(n40), .IN3(data3[12]), .IN4(n39), .Q(n27)
         );
  AO221X1 U31 ( .IN1(data1[11]), .IN2(n43), .IN3(data0[11]), .IN4(n42), .IN5(
        n26), .Q(data_o[11]) );
  AO22X1 U32 ( .IN1(data2[11]), .IN2(n40), .IN3(data3[11]), .IN4(n39), .Q(n26)
         );
  AO221X1 U33 ( .IN1(data1[10]), .IN2(n43), .IN3(data0[10]), .IN4(n42), .IN5(
        n25), .Q(data_o[10]) );
  AO22X1 U34 ( .IN1(data2[10]), .IN2(n40), .IN3(data3[10]), .IN4(n39), .Q(n25)
         );
  AO221X1 U35 ( .IN1(data1[0]), .IN2(n43), .IN3(data0[0]), .IN4(n42), .IN5(n24), .Q(data_o[0]) );
  AO22X1 U36 ( .IN1(data2[0]), .IN2(n40), .IN3(data3[0]), .IN4(n39), .Q(n24)
         );
  INVX0 U2 ( .INP(select2), .ZN(n1) );
  NOR4X0 U3 ( .IN1(n1), .IN2(select0), .IN3(select1), .IN4(select3), .QN(n40)
         );
  AND4X1 U4 ( .IN1(select3), .IN2(n3), .IN3(n2), .IN4(n1), .Q(n39) );
  INVX0 U37 ( .INP(select0), .ZN(n3) );
  INVX0 U38 ( .INP(select1), .ZN(n2) );
  NOR4X0 U39 ( .IN1(n3), .IN2(select1), .IN3(select2), .IN4(select3), .QN(n42)
         );
  NOR4X0 U40 ( .IN1(n2), .IN2(select0), .IN3(select2), .IN4(select3), .QN(n43)
         );
endmodule


module mux4_1_10 ( data0, data1, data2, data3, select0, select1, select2, 
        select3, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  input [15:0] data3;
  output [15:0] data_o;
  input select0, select1, select2, select3;
  wire   n1, n2, n3, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43;

  AO221X1 U5 ( .IN1(data1[9]), .IN2(n43), .IN3(data0[9]), .IN4(n42), .IN5(n41), 
        .Q(data_o[9]) );
  AO22X1 U6 ( .IN1(data2[9]), .IN2(n40), .IN3(data3[9]), .IN4(n39), .Q(n41) );
  AO221X1 U7 ( .IN1(data1[8]), .IN2(n43), .IN3(data0[8]), .IN4(n42), .IN5(n38), 
        .Q(data_o[8]) );
  AO22X1 U8 ( .IN1(data2[8]), .IN2(n40), .IN3(data3[8]), .IN4(n39), .Q(n38) );
  AO221X1 U9 ( .IN1(data1[7]), .IN2(n43), .IN3(data0[7]), .IN4(n42), .IN5(n37), 
        .Q(data_o[7]) );
  AO22X1 U10 ( .IN1(data2[7]), .IN2(n40), .IN3(data3[7]), .IN4(n39), .Q(n37)
         );
  AO221X1 U11 ( .IN1(data1[6]), .IN2(n43), .IN3(data0[6]), .IN4(n42), .IN5(n36), .Q(data_o[6]) );
  AO22X1 U12 ( .IN1(data2[6]), .IN2(n40), .IN3(data3[6]), .IN4(n39), .Q(n36)
         );
  AO221X1 U13 ( .IN1(data1[5]), .IN2(n43), .IN3(data0[5]), .IN4(n42), .IN5(n35), .Q(data_o[5]) );
  AO22X1 U14 ( .IN1(data2[5]), .IN2(n40), .IN3(data3[5]), .IN4(n39), .Q(n35)
         );
  AO221X1 U15 ( .IN1(data1[4]), .IN2(n43), .IN3(data0[4]), .IN4(n42), .IN5(n34), .Q(data_o[4]) );
  AO22X1 U16 ( .IN1(data2[4]), .IN2(n40), .IN3(data3[4]), .IN4(n39), .Q(n34)
         );
  AO221X1 U17 ( .IN1(data1[3]), .IN2(n43), .IN3(data0[3]), .IN4(n42), .IN5(n33), .Q(data_o[3]) );
  AO22X1 U18 ( .IN1(data2[3]), .IN2(n40), .IN3(data3[3]), .IN4(n39), .Q(n33)
         );
  AO221X1 U19 ( .IN1(data1[2]), .IN2(n43), .IN3(data0[2]), .IN4(n42), .IN5(n32), .Q(data_o[2]) );
  AO22X1 U20 ( .IN1(data2[2]), .IN2(n40), .IN3(data3[2]), .IN4(n39), .Q(n32)
         );
  AO221X1 U21 ( .IN1(data1[1]), .IN2(n43), .IN3(data0[1]), .IN4(n42), .IN5(n31), .Q(data_o[1]) );
  AO22X1 U22 ( .IN1(data2[1]), .IN2(n40), .IN3(data3[1]), .IN4(n39), .Q(n31)
         );
  AO221X1 U23 ( .IN1(data1[15]), .IN2(n43), .IN3(data0[15]), .IN4(n42), .IN5(
        n30), .Q(data_o[15]) );
  AO22X1 U24 ( .IN1(data2[15]), .IN2(n40), .IN3(data3[15]), .IN4(n39), .Q(n30)
         );
  AO221X1 U25 ( .IN1(data1[14]), .IN2(n43), .IN3(data0[14]), .IN4(n42), .IN5(
        n29), .Q(data_o[14]) );
  AO22X1 U26 ( .IN1(data2[14]), .IN2(n40), .IN3(data3[14]), .IN4(n39), .Q(n29)
         );
  AO221X1 U27 ( .IN1(data1[13]), .IN2(n43), .IN3(data0[13]), .IN4(n42), .IN5(
        n28), .Q(data_o[13]) );
  AO22X1 U28 ( .IN1(data2[13]), .IN2(n40), .IN3(data3[13]), .IN4(n39), .Q(n28)
         );
  AO221X1 U29 ( .IN1(data1[12]), .IN2(n43), .IN3(data0[12]), .IN4(n42), .IN5(
        n27), .Q(data_o[12]) );
  AO22X1 U30 ( .IN1(data2[12]), .IN2(n40), .IN3(data3[12]), .IN4(n39), .Q(n27)
         );
  AO221X1 U31 ( .IN1(data1[11]), .IN2(n43), .IN3(data0[11]), .IN4(n42), .IN5(
        n26), .Q(data_o[11]) );
  AO22X1 U32 ( .IN1(data2[11]), .IN2(n40), .IN3(data3[11]), .IN4(n39), .Q(n26)
         );
  AO221X1 U33 ( .IN1(data1[10]), .IN2(n43), .IN3(data0[10]), .IN4(n42), .IN5(
        n25), .Q(data_o[10]) );
  AO22X1 U34 ( .IN1(data2[10]), .IN2(n40), .IN3(data3[10]), .IN4(n39), .Q(n25)
         );
  AO221X1 U35 ( .IN1(data1[0]), .IN2(n43), .IN3(data0[0]), .IN4(n42), .IN5(n24), .Q(data_o[0]) );
  AO22X1 U36 ( .IN1(data2[0]), .IN2(n40), .IN3(data3[0]), .IN4(n39), .Q(n24)
         );
  INVX0 U2 ( .INP(select2), .ZN(n1) );
  NOR4X0 U3 ( .IN1(n1), .IN2(select0), .IN3(select1), .IN4(select3), .QN(n40)
         );
  AND4X1 U4 ( .IN1(select3), .IN2(n3), .IN3(n2), .IN4(n1), .Q(n39) );
  INVX0 U37 ( .INP(select0), .ZN(n3) );
  INVX0 U38 ( .INP(select1), .ZN(n2) );
  NOR4X0 U39 ( .IN1(n3), .IN2(select1), .IN3(select2), .IN4(select3), .QN(n42)
         );
  NOR4X0 U40 ( .IN1(n2), .IN2(select0), .IN3(select2), .IN4(select3), .QN(n43)
         );
endmodule


module mux4_1_9 ( data0, data1, data2, data3, select0, select1, select2, 
        select3, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  input [15:0] data3;
  output [15:0] data_o;
  input select0, select1, select2, select3;
  wire   n1, n2, n3, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43;

  AO221X1 U5 ( .IN1(data1[9]), .IN2(n43), .IN3(data0[9]), .IN4(n42), .IN5(n41), 
        .Q(data_o[9]) );
  AO22X1 U6 ( .IN1(data2[9]), .IN2(n40), .IN3(data3[9]), .IN4(n39), .Q(n41) );
  AO221X1 U7 ( .IN1(data1[8]), .IN2(n43), .IN3(data0[8]), .IN4(n42), .IN5(n38), 
        .Q(data_o[8]) );
  AO22X1 U8 ( .IN1(data2[8]), .IN2(n40), .IN3(data3[8]), .IN4(n39), .Q(n38) );
  AO221X1 U9 ( .IN1(data1[7]), .IN2(n43), .IN3(data0[7]), .IN4(n42), .IN5(n37), 
        .Q(data_o[7]) );
  AO22X1 U10 ( .IN1(data2[7]), .IN2(n40), .IN3(data3[7]), .IN4(n39), .Q(n37)
         );
  AO221X1 U11 ( .IN1(data1[6]), .IN2(n43), .IN3(data0[6]), .IN4(n42), .IN5(n36), .Q(data_o[6]) );
  AO22X1 U12 ( .IN1(data2[6]), .IN2(n40), .IN3(data3[6]), .IN4(n39), .Q(n36)
         );
  AO221X1 U13 ( .IN1(data1[5]), .IN2(n43), .IN3(data0[5]), .IN4(n42), .IN5(n35), .Q(data_o[5]) );
  AO22X1 U14 ( .IN1(data2[5]), .IN2(n40), .IN3(data3[5]), .IN4(n39), .Q(n35)
         );
  AO221X1 U15 ( .IN1(data1[4]), .IN2(n43), .IN3(data0[4]), .IN4(n42), .IN5(n34), .Q(data_o[4]) );
  AO22X1 U16 ( .IN1(data2[4]), .IN2(n40), .IN3(data3[4]), .IN4(n39), .Q(n34)
         );
  AO221X1 U17 ( .IN1(data1[3]), .IN2(n43), .IN3(data0[3]), .IN4(n42), .IN5(n33), .Q(data_o[3]) );
  AO22X1 U18 ( .IN1(data2[3]), .IN2(n40), .IN3(data3[3]), .IN4(n39), .Q(n33)
         );
  AO221X1 U19 ( .IN1(data1[2]), .IN2(n43), .IN3(data0[2]), .IN4(n42), .IN5(n32), .Q(data_o[2]) );
  AO22X1 U20 ( .IN1(data2[2]), .IN2(n40), .IN3(data3[2]), .IN4(n39), .Q(n32)
         );
  AO221X1 U21 ( .IN1(data1[1]), .IN2(n43), .IN3(data0[1]), .IN4(n42), .IN5(n31), .Q(data_o[1]) );
  AO22X1 U22 ( .IN1(data2[1]), .IN2(n40), .IN3(data3[1]), .IN4(n39), .Q(n31)
         );
  AO221X1 U23 ( .IN1(data1[15]), .IN2(n43), .IN3(data0[15]), .IN4(n42), .IN5(
        n30), .Q(data_o[15]) );
  AO22X1 U24 ( .IN1(data2[15]), .IN2(n40), .IN3(data3[15]), .IN4(n39), .Q(n30)
         );
  AO221X1 U25 ( .IN1(data1[14]), .IN2(n43), .IN3(data0[14]), .IN4(n42), .IN5(
        n29), .Q(data_o[14]) );
  AO22X1 U26 ( .IN1(data2[14]), .IN2(n40), .IN3(data3[14]), .IN4(n39), .Q(n29)
         );
  AO221X1 U27 ( .IN1(data1[13]), .IN2(n43), .IN3(data0[13]), .IN4(n42), .IN5(
        n28), .Q(data_o[13]) );
  AO22X1 U28 ( .IN1(data2[13]), .IN2(n40), .IN3(data3[13]), .IN4(n39), .Q(n28)
         );
  AO221X1 U29 ( .IN1(data1[12]), .IN2(n43), .IN3(data0[12]), .IN4(n42), .IN5(
        n27), .Q(data_o[12]) );
  AO22X1 U30 ( .IN1(data2[12]), .IN2(n40), .IN3(data3[12]), .IN4(n39), .Q(n27)
         );
  AO221X1 U31 ( .IN1(data1[11]), .IN2(n43), .IN3(data0[11]), .IN4(n42), .IN5(
        n26), .Q(data_o[11]) );
  AO22X1 U32 ( .IN1(data2[11]), .IN2(n40), .IN3(data3[11]), .IN4(n39), .Q(n26)
         );
  AO221X1 U33 ( .IN1(data1[10]), .IN2(n43), .IN3(data0[10]), .IN4(n42), .IN5(
        n25), .Q(data_o[10]) );
  AO22X1 U34 ( .IN1(data2[10]), .IN2(n40), .IN3(data3[10]), .IN4(n39), .Q(n25)
         );
  AO221X1 U35 ( .IN1(data1[0]), .IN2(n43), .IN3(data0[0]), .IN4(n42), .IN5(n24), .Q(data_o[0]) );
  AO22X1 U36 ( .IN1(data2[0]), .IN2(n40), .IN3(data3[0]), .IN4(n39), .Q(n24)
         );
  INVX0 U2 ( .INP(select2), .ZN(n1) );
  NOR4X0 U3 ( .IN1(n1), .IN2(select0), .IN3(select1), .IN4(select3), .QN(n40)
         );
  AND4X1 U4 ( .IN1(select3), .IN2(n3), .IN3(n2), .IN4(n1), .Q(n39) );
  INVX0 U37 ( .INP(select0), .ZN(n3) );
  INVX0 U38 ( .INP(select1), .ZN(n2) );
  NOR4X0 U39 ( .IN1(n3), .IN2(select1), .IN3(select2), .IN4(select3), .QN(n42)
         );
  NOR4X0 U40 ( .IN1(n2), .IN2(select0), .IN3(select2), .IN4(select3), .QN(n43)
         );
endmodule



    module node5_NODE_X1_NODE_Y1I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__I_node_2_node_interface__I_node_3_node_interface__ ( 
        \clk.clk , \reset.reset , \local_node.clk , 
        \local_node.buffer_full_in , \local_node.buffer_full_out , 
        \local_node.receiving_data , \local_node.sending_data , 
        \local_node.data_in , \local_node.data_out , \node_0.clk , 
        \node_0.buffer_full_in , \node_0.buffer_full_out , 
        \node_0.receiving_data , \node_0.sending_data , \node_0.data_in , 
        \node_0.data_out , \node_1.clk , \node_1.buffer_full_in , 
        \node_1.buffer_full_out , \node_1.receiving_data , 
        \node_1.sending_data , \node_1.data_in , \node_1.data_out , 
        \node_2.clk , \node_2.buffer_full_in , \node_2.buffer_full_out , 
        \node_2.receiving_data , \node_2.sending_data , \node_2.data_in , 
        \node_2.data_out , \node_3.clk , \node_3.buffer_full_in , 
        \node_3.buffer_full_out , \node_3.receiving_data , 
        \node_3.sending_data , \node_3.data_in , \node_3.data_out  );
  input [15:0] \local_node.data_in ;
  output [15:0] \local_node.data_out ;
  input [15:0] \node_0.data_in ;
  output [15:0] \node_0.data_out ;
  input [15:0] \node_1.data_in ;
  output [15:0] \node_1.data_out ;
  input [15:0] \node_2.data_in ;
  output [15:0] \node_2.data_out ;
  input [15:0] \node_3.data_in ;
  output [15:0] \node_3.data_out ;
  input \clk.clk , \reset.reset , \local_node.buffer_full_in ,
         \local_node.receiving_data , \node_0.buffer_full_in ,
         \node_0.receiving_data , \node_1.buffer_full_in ,
         \node_1.receiving_data , \node_2.buffer_full_in ,
         \node_2.receiving_data , \node_3.buffer_full_in ,
         \node_3.receiving_data ;
  output \local_node.buffer_full_out , \local_node.sending_data ,
         \node_0.buffer_full_out , \node_0.sending_data ,
         \node_1.buffer_full_out , \node_1.sending_data ,
         \node_2.buffer_full_out , \node_2.sending_data ,
         \node_3.buffer_full_out , \node_3.sending_data ;
  inout \local_node.clk ,  \node_0.clk ,  \node_1.clk ,  \node_2.clk , 
     \node_3.clk ;
  wire   \buffer_out[4][15] , \buffer_out[4][14] , \buffer_out[4][13] ,
         \buffer_out[4][12] , \buffer_out[4][11] , \buffer_out[4][10] ,
         \buffer_out[4][9] , \buffer_out[4][8] , \buffer_out[4][7] ,
         \buffer_out[4][6] , \buffer_out[4][5] , \buffer_out[4][4] ,
         \buffer_out[4][3] , \buffer_out[4][2] , \buffer_out[4][1] ,
         \buffer_out[4][0] , \buffer_out[3][15] , \buffer_out[3][14] ,
         \buffer_out[3][13] , \buffer_out[3][12] , \buffer_out[3][11] ,
         \buffer_out[3][10] , \buffer_out[3][9] , \buffer_out[3][8] ,
         \buffer_out[3][7] , \buffer_out[3][6] , \buffer_out[3][5] ,
         \buffer_out[3][4] , \buffer_out[3][3] , \buffer_out[3][2] ,
         \buffer_out[3][1] , \buffer_out[3][0] , \buffer_out[2][15] ,
         \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] ,
         \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] ,
         \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] ,
         \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] ,
         \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] ,
         \buffer_out[1][15] , \buffer_out[1][14] , \buffer_out[1][13] ,
         \buffer_out[1][12] , \buffer_out[1][11] , \buffer_out[1][10] ,
         \buffer_out[1][9] , \buffer_out[1][8] , \buffer_out[1][7] ,
         \buffer_out[1][6] , \buffer_out[1][5] , \buffer_out[1][4] ,
         \buffer_out[1][3] , \buffer_out[1][2] , \buffer_out[1][1] ,
         \buffer_out[1][0] , \buffer_out[0][15] , \buffer_out[0][14] ,
         \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] ,
         \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] ,
         \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] ,
         \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] ,
         \buffer_out[0][1] , \buffer_out[0][0] , \next_buffer_out[4][15] ,
         \next_buffer_out[4][14] , \next_buffer_out[4][13] ,
         \next_buffer_out[4][12] , \next_buffer_out[4][11] ,
         \next_buffer_out[4][10] , \next_buffer_out[4][9] ,
         \next_buffer_out[4][8] , \next_buffer_out[4][7] ,
         \next_buffer_out[4][6] , \next_buffer_out[4][5] ,
         \next_buffer_out[4][4] , \next_buffer_out[4][3] ,
         \next_buffer_out[4][2] , \next_buffer_out[4][1] ,
         \next_buffer_out[4][0] , \next_buffer_out[3][15] ,
         \next_buffer_out[3][14] , \next_buffer_out[3][13] ,
         \next_buffer_out[3][12] , \next_buffer_out[3][11] ,
         \next_buffer_out[3][10] , \next_buffer_out[3][9] ,
         \next_buffer_out[3][8] , \next_buffer_out[3][7] ,
         \next_buffer_out[3][6] , \next_buffer_out[3][5] ,
         \next_buffer_out[3][4] , \next_buffer_out[3][3] ,
         \next_buffer_out[3][2] , \next_buffer_out[3][1] ,
         \next_buffer_out[3][0] , \next_buffer_out[2][15] ,
         \next_buffer_out[2][14] , \next_buffer_out[2][13] ,
         \next_buffer_out[2][12] , \next_buffer_out[2][11] ,
         \next_buffer_out[2][10] , \next_buffer_out[2][9] ,
         \next_buffer_out[2][8] , \next_buffer_out[2][7] ,
         \next_buffer_out[2][6] , \next_buffer_out[2][5] ,
         \next_buffer_out[2][4] , \next_buffer_out[2][3] ,
         \next_buffer_out[2][2] , \next_buffer_out[2][1] ,
         \next_buffer_out[2][0] , \next_buffer_out[1][15] ,
         \next_buffer_out[1][14] , \next_buffer_out[1][13] ,
         \next_buffer_out[1][12] , \next_buffer_out[1][11] ,
         \next_buffer_out[1][10] , \next_buffer_out[1][9] ,
         \next_buffer_out[1][8] , \next_buffer_out[1][7] ,
         \next_buffer_out[1][6] , \next_buffer_out[1][5] ,
         \next_buffer_out[1][4] , \next_buffer_out[1][3] ,
         \next_buffer_out[1][2] , \next_buffer_out[1][1] ,
         \next_buffer_out[1][0] , \next_buffer_out[0][15] ,
         \next_buffer_out[0][14] , \next_buffer_out[0][13] ,
         \next_buffer_out[0][12] , \next_buffer_out[0][11] ,
         \next_buffer_out[0][10] , \next_buffer_out[0][9] ,
         \next_buffer_out[0][8] , \next_buffer_out[0][7] ,
         \next_buffer_out[0][6] , \next_buffer_out[0][5] ,
         \next_buffer_out[0][4] , \next_buffer_out[0][3] ,
         \next_buffer_out[0][2] , \next_buffer_out[0][1] ,
         \next_buffer_out[0][0] ;
  wire   [4:0] buffer_full_in;
  wire   [4:0] receiving_data;
  wire   [4:0] pop_v;
  wire   [4:0] data_valid;
  wire   [4:0] next_data_valid;
  wire   [1:0] grant_0;
  wire   [1:0] grant_1;
  wire   [3:0] grant_2;
  wire   [3:0] grant_3;
  wire   [3:0] grant_4;
  tri   \local_node.buffer_full_in ;
  tri   \local_node.buffer_full_out ;
  tri   \local_node.receiving_data ;
  tri   \local_node.sending_data ;
  tri   [15:0] \local_node.data_in ;
  tri   [15:0] \local_node.data_out ;

  converter_in_I_n_node_interface_dut__7 c0 ( .\n.buffer_full_in (
        \node_0.buffer_full_in ), .\n.receiving_data (\node_0.receiving_data ), 
        .\n.data_in (\node_0.data_in ), .\n.buffer_full_out (
        \node_0.buffer_full_out ), .\n.sending_data (\node_0.sending_data ), 
        .\n.data_out (\node_0.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_out_I_n_node_interface_dut_ c1 ( .\n.buffer_full_in (
        \node_1.buffer_full_in ), .\n.receiving_data (\node_1.receiving_data ), 
        .\n.data_in (\node_1.data_in ), .\n.buffer_full_out (
        \node_1.buffer_full_out ), .\n.sending_data (\node_1.sending_data ), 
        .\n.data_out (\node_1.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_in_I_n_node_interface_dut__6 c2 ( .\n.buffer_full_in (
        \node_2.buffer_full_in ), .\n.receiving_data (\node_2.receiving_data ), 
        .\n.data_in (\node_2.data_in ), .\n.buffer_full_out (
        \node_2.buffer_full_out ), .\n.sending_data (\node_2.sending_data ), 
        .\n.data_out (\node_2.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_out_I_n_node_interface_dut_ c3 ( .\n.buffer_full_in (
        \node_3.buffer_full_in ), .\n.receiving_data (\node_3.receiving_data ), 
        .\n.data_in (\node_3.data_in ), .\n.buffer_full_out (
        \node_3.buffer_full_out ), .\n.sending_data (\node_3.sending_data ), 
        .\n.data_out (\node_3.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_out_I_n_node_interface_dut_ c4 ( .\n.buffer_full_in (
        \local_node.buffer_full_in ), .\n.receiving_data (
        \local_node.receiving_data ), .\n.data_in (\local_node.data_in ), 
        .\n.buffer_full_out (\local_node.buffer_full_out ), .\n.sending_data (
        \local_node.sending_data ), .\n.data_out (\local_node.data_out ), 
        .buffer_full_in(1'b0), .receiving_data(1'b0), .data_in({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  fifo_kev_19 \genblk1[0].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[0]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[0]), .data_out({\buffer_out[0][15] , 
        \buffer_out[0][14] , \buffer_out[0][13] , \buffer_out[0][12] , 
        \buffer_out[0][11] , \buffer_out[0][10] , \buffer_out[0][9] , 
        \buffer_out[0][8] , \buffer_out[0][7] , \buffer_out[0][6] , 
        \buffer_out[0][5] , \buffer_out[0][4] , \buffer_out[0][3] , 
        \buffer_out[0][2] , \buffer_out[0][1] , \buffer_out[0][0] }), 
        .next_data_out({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] , 
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .next_data_valid(
        next_data_valid[0]) );
  address_counter_19 \genblk1[0].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] }), 
        .buffer_data_valid(next_data_valid[0]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .buffer_pop(
        pop_v[0]), .receiving_data(1'b0) );
  fifo_kev_18 \genblk1[1].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[1]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[1]), .data_out({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), 
        .next_data_out({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] , 
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .next_data_valid(
        next_data_valid[1]) );
  address_counter_18 \genblk1[1].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] }), 
        .buffer_data_valid(next_data_valid[1]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .buffer_pop(
        pop_v[1]), .receiving_data(1'b0) );
  fifo_kev_17 \genblk1[2].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[2]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[2]), .data_out({\buffer_out[2][15] , 
        \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] , 
        \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] , 
        \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] , 
        \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] , 
        \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] }), 
        .next_data_out({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] , 
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .next_data_valid(
        next_data_valid[2]) );
  address_counter_17 \genblk1[2].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] }), 
        .buffer_data_valid(next_data_valid[2]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .buffer_pop(
        pop_v[2]), .receiving_data(1'b0) );
  fifo_kev_16 \genblk1[3].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[3]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[3]), .data_out({\buffer_out[3][15] , 
        \buffer_out[3][14] , \buffer_out[3][13] , \buffer_out[3][12] , 
        \buffer_out[3][11] , \buffer_out[3][10] , \buffer_out[3][9] , 
        \buffer_out[3][8] , \buffer_out[3][7] , \buffer_out[3][6] , 
        \buffer_out[3][5] , \buffer_out[3][4] , \buffer_out[3][3] , 
        \buffer_out[3][2] , \buffer_out[3][1] , \buffer_out[3][0] }), 
        .next_data_out({\next_buffer_out[3][15] , \next_buffer_out[3][14] , 
        \next_buffer_out[3][13] , \next_buffer_out[3][12] , 
        \next_buffer_out[3][11] , \next_buffer_out[3][10] , 
        \next_buffer_out[3][9] , \next_buffer_out[3][8] , 
        \next_buffer_out[3][7] , \next_buffer_out[3][6] , 
        \next_buffer_out[3][5] , \next_buffer_out[3][4] , 
        \next_buffer_out[3][3] , \next_buffer_out[3][2] , 
        \next_buffer_out[3][1] , \next_buffer_out[3][0] }), .next_data_valid(
        next_data_valid[3]) );
  address_counter_16 \genblk1[3].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[3][15] , \next_buffer_out[3][14] , 
        \next_buffer_out[3][13] , \next_buffer_out[3][12] , 
        \next_buffer_out[3][11] , \next_buffer_out[3][10] , 
        \next_buffer_out[3][9] , \next_buffer_out[3][8] }), 
        .buffer_data_valid(next_data_valid[3]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[3][7] , \next_buffer_out[3][6] , 
        \next_buffer_out[3][5] , \next_buffer_out[3][4] , 
        \next_buffer_out[3][3] , \next_buffer_out[3][2] , 
        \next_buffer_out[3][1] , \next_buffer_out[3][0] }), .buffer_pop(
        pop_v[3]), .receiving_data(1'b0) );
  fifo_kev_15 \genblk1[4].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[4]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[4]), .data_out({\buffer_out[4][15] , 
        \buffer_out[4][14] , \buffer_out[4][13] , \buffer_out[4][12] , 
        \buffer_out[4][11] , \buffer_out[4][10] , \buffer_out[4][9] , 
        \buffer_out[4][8] , \buffer_out[4][7] , \buffer_out[4][6] , 
        \buffer_out[4][5] , \buffer_out[4][4] , \buffer_out[4][3] , 
        \buffer_out[4][2] , \buffer_out[4][1] , \buffer_out[4][0] }), 
        .next_data_out({\next_buffer_out[4][15] , \next_buffer_out[4][14] , 
        \next_buffer_out[4][13] , \next_buffer_out[4][12] , 
        \next_buffer_out[4][11] , \next_buffer_out[4][10] , 
        \next_buffer_out[4][9] , \next_buffer_out[4][8] , 
        \next_buffer_out[4][7] , \next_buffer_out[4][6] , 
        \next_buffer_out[4][5] , \next_buffer_out[4][4] , 
        \next_buffer_out[4][3] , \next_buffer_out[4][2] , 
        \next_buffer_out[4][1] , \next_buffer_out[4][0] }), .next_data_valid(
        next_data_valid[4]) );
  address_counter_15 \genblk1[4].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[4][15] , \next_buffer_out[4][14] , 
        \next_buffer_out[4][13] , \next_buffer_out[4][12] , 
        \next_buffer_out[4][11] , \next_buffer_out[4][10] , 
        \next_buffer_out[4][9] , \next_buffer_out[4][8] }), 
        .buffer_data_valid(next_data_valid[4]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[4][7] , \next_buffer_out[4][6] , 
        \next_buffer_out[4][5] , \next_buffer_out[4][4] , 
        \next_buffer_out[4][3] , \next_buffer_out[4][2] , 
        \next_buffer_out[4][1] , \next_buffer_out[4][0] }), .buffer_pop(
        pop_v[4]), .receiving_data(1'b0) );
  controller5_3 ctrl5 ( .clk(\clk.clk ), .rst(\reset.reset ), .packet_addr({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .local_addr({1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 
        1'b0, 1'b0, 1'b1}), .packet_valid(data_valid), .buffer_full_in({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .grant_0(grant_0), .grant_1(grant_1), 
        .grant_2(grant_2), .grant_3(grant_3), .grant_4(grant_4), .pop_v(pop_v)
         );
  mux2_1_7 mux_n ( .data0({\buffer_out[1][15] , \buffer_out[1][14] , 
        \buffer_out[1][13] , \buffer_out[1][12] , \buffer_out[1][11] , 
        \buffer_out[1][10] , \buffer_out[1][9] , \buffer_out[1][8] , 
        \buffer_out[1][7] , \buffer_out[1][6] , \buffer_out[1][5] , 
        \buffer_out[1][4] , \buffer_out[1][3] , \buffer_out[1][2] , 
        \buffer_out[1][1] , \buffer_out[1][0] }), .data1({\buffer_out[4][15] , 
        \buffer_out[4][14] , \buffer_out[4][13] , \buffer_out[4][12] , 
        \buffer_out[4][11] , \buffer_out[4][10] , \buffer_out[4][9] , 
        \buffer_out[4][8] , \buffer_out[4][7] , \buffer_out[4][6] , 
        \buffer_out[4][5] , \buffer_out[4][4] , \buffer_out[4][3] , 
        \buffer_out[4][2] , \buffer_out[4][1] , \buffer_out[4][0] }), 
        .select0(grant_0[0]), .select1(grant_0[1]) );
  mux2_1_6 mux_s ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[4][15] , 
        \buffer_out[4][14] , \buffer_out[4][13] , \buffer_out[4][12] , 
        \buffer_out[4][11] , \buffer_out[4][10] , \buffer_out[4][9] , 
        \buffer_out[4][8] , \buffer_out[4][7] , \buffer_out[4][6] , 
        \buffer_out[4][5] , \buffer_out[4][4] , \buffer_out[4][3] , 
        \buffer_out[4][2] , \buffer_out[4][1] , \buffer_out[4][0] }), 
        .select0(grant_1[0]), .select1(grant_1[1]) );
  mux4_1_11 mux_e ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[3][15] , \buffer_out[3][14] , \buffer_out[3][13] , 
        \buffer_out[3][12] , \buffer_out[3][11] , \buffer_out[3][10] , 
        \buffer_out[3][9] , \buffer_out[3][8] , \buffer_out[3][7] , 
        \buffer_out[3][6] , \buffer_out[3][5] , \buffer_out[3][4] , 
        \buffer_out[3][3] , \buffer_out[3][2] , \buffer_out[3][1] , 
        \buffer_out[3][0] }), .data3({\buffer_out[4][15] , \buffer_out[4][14] , 
        \buffer_out[4][13] , \buffer_out[4][12] , \buffer_out[4][11] , 
        \buffer_out[4][10] , \buffer_out[4][9] , \buffer_out[4][8] , 
        \buffer_out[4][7] , \buffer_out[4][6] , \buffer_out[4][5] , 
        \buffer_out[4][4] , \buffer_out[4][3] , \buffer_out[4][2] , 
        \buffer_out[4][1] , \buffer_out[4][0] }), .select0(grant_2[0]), 
        .select1(grant_2[1]), .select2(grant_2[2]), .select3(grant_2[3]) );
  mux4_1_10 mux_w ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[2][15] , \buffer_out[2][14] , \buffer_out[2][13] , 
        \buffer_out[2][12] , \buffer_out[2][11] , \buffer_out[2][10] , 
        \buffer_out[2][9] , \buffer_out[2][8] , \buffer_out[2][7] , 
        \buffer_out[2][6] , \buffer_out[2][5] , \buffer_out[2][4] , 
        \buffer_out[2][3] , \buffer_out[2][2] , \buffer_out[2][1] , 
        \buffer_out[2][0] }), .data3({\buffer_out[4][15] , \buffer_out[4][14] , 
        \buffer_out[4][13] , \buffer_out[4][12] , \buffer_out[4][11] , 
        \buffer_out[4][10] , \buffer_out[4][9] , \buffer_out[4][8] , 
        \buffer_out[4][7] , \buffer_out[4][6] , \buffer_out[4][5] , 
        \buffer_out[4][4] , \buffer_out[4][3] , \buffer_out[4][2] , 
        \buffer_out[4][1] , \buffer_out[4][0] }), .select0(grant_3[0]), 
        .select1(grant_3[1]), .select2(grant_3[2]), .select3(grant_3[3]) );
  mux4_1_9 mux_l ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[2][15] , \buffer_out[2][14] , \buffer_out[2][13] , 
        \buffer_out[2][12] , \buffer_out[2][11] , \buffer_out[2][10] , 
        \buffer_out[2][9] , \buffer_out[2][8] , \buffer_out[2][7] , 
        \buffer_out[2][6] , \buffer_out[2][5] , \buffer_out[2][4] , 
        \buffer_out[2][3] , \buffer_out[2][2] , \buffer_out[2][1] , 
        \buffer_out[2][0] }), .data3({\buffer_out[3][15] , \buffer_out[3][14] , 
        \buffer_out[3][13] , \buffer_out[3][12] , \buffer_out[3][11] , 
        \buffer_out[3][10] , \buffer_out[3][9] , \buffer_out[3][8] , 
        \buffer_out[3][7] , \buffer_out[3][6] , \buffer_out[3][5] , 
        \buffer_out[3][4] , \buffer_out[3][3] , \buffer_out[3][2] , 
        \buffer_out[3][1] , \buffer_out[3][0] }), .select0(grant_4[0]), 
        .select1(grant_4[1]), .select2(grant_4[2]), .select3(grant_4[3]) );
endmodule


module converter_in_I_n_node_interface_dut__5 ( \n.buffer_full_in , 
        \n.receiving_data , \n.data_in , \n.buffer_full_out , \n.sending_data , 
        \n.data_out , buffer_full_out, sending_data, data_out, buffer_full_in, 
        receiving_data, data_in );
  input [15:0] \n.data_in ;
  output [15:0] \n.data_out ;
  output [15:0] data_out;
  input [15:0] data_in;
  input \n.buffer_full_in , \n.receiving_data , buffer_full_in, receiving_data;
  output \n.buffer_full_out , \n.sending_data , buffer_full_out, sending_data;
  wire   \n.buffer_full_in , \n.receiving_data , buffer_full_in,
         receiving_data;
  assign buffer_full_out = \n.buffer_full_in ;
  assign sending_data = \n.receiving_data ;
  assign data_out[15] = \n.data_in  [15];
  assign data_out[14] = \n.data_in  [14];
  assign data_out[13] = \n.data_in  [13];
  assign data_out[12] = \n.data_in  [12];
  assign data_out[11] = \n.data_in  [11];
  assign data_out[10] = \n.data_in  [10];
  assign data_out[9] = \n.data_in  [9];
  assign data_out[8] = \n.data_in  [8];
  assign data_out[7] = \n.data_in  [7];
  assign data_out[6] = \n.data_in  [6];
  assign data_out[5] = \n.data_in  [5];
  assign data_out[4] = \n.data_in  [4];
  assign data_out[3] = \n.data_in  [3];
  assign data_out[2] = \n.data_in  [2];
  assign data_out[1] = \n.data_in  [1];
  assign data_out[0] = \n.data_in  [0];
  assign \n.buffer_full_out  = buffer_full_in;
  assign \n.sending_data  = receiving_data;
  assign \n.data_out  [15] = data_in[15];
  assign \n.data_out  [14] = data_in[14];
  assign \n.data_out  [13] = data_in[13];
  assign \n.data_out  [12] = data_in[12];
  assign \n.data_out  [11] = data_in[11];
  assign \n.data_out  [10] = data_in[10];
  assign \n.data_out  [9] = data_in[9];
  assign \n.data_out  [8] = data_in[8];
  assign \n.data_out  [7] = data_in[7];
  assign \n.data_out  [6] = data_in[6];
  assign \n.data_out  [5] = data_in[5];
  assign \n.data_out  [4] = data_in[4];
  assign \n.data_out  [3] = data_in[3];
  assign \n.data_out  [2] = data_in[2];
  assign \n.data_out  [1] = data_in[1];
  assign \n.data_out  [0] = data_in[0];

endmodule


module converter_in_I_n_node_interface_dut__4 ( \n.buffer_full_in , 
        \n.receiving_data , \n.data_in , \n.buffer_full_out , \n.sending_data , 
        \n.data_out , buffer_full_out, sending_data, data_out, buffer_full_in, 
        receiving_data, data_in );
  input [15:0] \n.data_in ;
  output [15:0] \n.data_out ;
  output [15:0] data_out;
  input [15:0] data_in;
  input \n.buffer_full_in , \n.receiving_data , buffer_full_in, receiving_data;
  output \n.buffer_full_out , \n.sending_data , buffer_full_out, sending_data;
  wire   \n.buffer_full_in , \n.receiving_data , buffer_full_in,
         receiving_data;
  assign buffer_full_out = \n.buffer_full_in ;
  assign sending_data = \n.receiving_data ;
  assign data_out[15] = \n.data_in  [15];
  assign data_out[14] = \n.data_in  [14];
  assign data_out[13] = \n.data_in  [13];
  assign data_out[12] = \n.data_in  [12];
  assign data_out[11] = \n.data_in  [11];
  assign data_out[10] = \n.data_in  [10];
  assign data_out[9] = \n.data_in  [9];
  assign data_out[8] = \n.data_in  [8];
  assign data_out[7] = \n.data_in  [7];
  assign data_out[6] = \n.data_in  [6];
  assign data_out[5] = \n.data_in  [5];
  assign data_out[4] = \n.data_in  [4];
  assign data_out[3] = \n.data_in  [3];
  assign data_out[2] = \n.data_in  [2];
  assign data_out[1] = \n.data_in  [1];
  assign data_out[0] = \n.data_in  [0];
  assign \n.buffer_full_out  = buffer_full_in;
  assign \n.sending_data  = receiving_data;
  assign \n.data_out  [15] = data_in[15];
  assign \n.data_out  [14] = data_in[14];
  assign \n.data_out  [13] = data_in[13];
  assign \n.data_out  [12] = data_in[12];
  assign \n.data_out  [11] = data_in[11];
  assign \n.data_out  [10] = data_in[10];
  assign \n.data_out  [9] = data_in[9];
  assign \n.data_out  [8] = data_in[8];
  assign \n.data_out  [7] = data_in[7];
  assign \n.data_out  [6] = data_in[6];
  assign \n.data_out  [5] = data_in[5];
  assign \n.data_out  [4] = data_in[4];
  assign \n.data_out  [3] = data_in[3];
  assign \n.data_out  [2] = data_in[2];
  assign \n.data_out  [1] = data_in[1];
  assign \n.data_out  [0] = data_in[0];

endmodule


module fifo_kev_14 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_29 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_14 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_29 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_28 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_14 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_28 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_14_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_14 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_14 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_14 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_14_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_13 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_27 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_13 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_27 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_26 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_13 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_26 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_13_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_13 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_13 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_13 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_13_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_12 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_25 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_12 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_25 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_24 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_12 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_24 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_12_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_12 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_12 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_12 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_12_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_11 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_23 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_11 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_23 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_22 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_11 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_22 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_11_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_11 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_11 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_11 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_11_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_10 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_21 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_10 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_21 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_20 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_10 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_20 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_10_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_10 ( clk, rst, interface_flit_length, 
        buffer_flit_length, buffer_data_valid, interface_flit_address, 
        buffer_flit_address, buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_10 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_10 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_10_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module flipflop_BITS2_5 ( clk, data_i, data_o );
  input [1:0] data_i;
  output [1:0] data_o;
  input clk;


  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS2_5 ( clk, enable_i, reset, data_i, data_o );
  input [1:0] data_i;
  input [1:0] data_o;
  input clk, enable_i, reset;
  wire   n10, n11, n1, n5, n7, n8, n9;
  wire   [1:0] write_data;

  AOI22X1 U5 ( .IN1(enable_i), .IN2(data_i[1]), .IN3(n10), .IN4(n1), .QN(n9)
         );
  AOI22X1 U6 ( .IN1(data_i[0]), .IN2(enable_i), .IN3(n11), .IN4(n1), .QN(n8)
         );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n9), .QN(write_data[1]) );
  NOR2X0 U4 ( .IN1(reset), .IN2(n8), .QN(write_data[0]) );
  AND2X1 U7 ( .IN1(data_o[1]), .IN2(n7), .Q(n10) );
  AND2X1 U8 ( .IN1(data_o[0]), .IN2(n5), .Q(n11) );
  flipflop_BITS2_5 FF ( .clk(clk), .data_i(write_data), .data_o({n7, n5}) );
endmodule


module flipflop_BITS1_23 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_23 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_23 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter2_5 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [1:0] request;
  output [1:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   tail_en, n1, n2;
  wire   [1:0] req_i;
  wire   [1:0] req_o;

  AND3X1 U10 ( .IN1(request[1]), .IN2(n1), .IN3(n2), .Q(grant[1]) );
  AND3X1 U11 ( .IN1(request[0]), .IN2(n2), .IN3(request[1]), .Q(tail_en) );
  INVX0 U6 ( .INP(request[0]), .ZN(n1) );
  NOR2X0 U7 ( .IN1(buffer_full_i), .IN2(n1), .QN(grant[0]) );
  INVX0 U8 ( .INP(buffer_full_i), .ZN(n2) );
  OA21X1 U9 ( .IN1(request[1]), .IN2(request[0]), .IN3(n2), .Q(grant_v_o) );
  register_BITS2_5 req_record ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i({1'b1, 1'b0}), .data_o({1'b0, 1'b0}) );
  register_BITS1_23 tail ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i(1'b1), .data_o(1'b0) );
endmodule


module flipflop_BITS2_4 ( clk, data_i, data_o );
  input [1:0] data_i;
  output [1:0] data_o;
  input clk;


  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS2_4 ( clk, enable_i, reset, data_i, data_o );
  input [1:0] data_i;
  input [1:0] data_o;
  input clk, enable_i, reset;
  wire   n10, n11, n1, n5, n7, n8, n9;
  wire   [1:0] write_data;

  AOI22X1 U5 ( .IN1(enable_i), .IN2(data_i[1]), .IN3(n10), .IN4(n1), .QN(n9)
         );
  AOI22X1 U6 ( .IN1(data_i[0]), .IN2(enable_i), .IN3(n11), .IN4(n1), .QN(n8)
         );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n9), .QN(write_data[1]) );
  NOR2X0 U4 ( .IN1(reset), .IN2(n8), .QN(write_data[0]) );
  AND2X1 U7 ( .IN1(data_o[1]), .IN2(n7), .Q(n10) );
  AND2X1 U8 ( .IN1(data_o[0]), .IN2(n5), .Q(n11) );
  flipflop_BITS2_4 FF ( .clk(clk), .data_i(write_data), .data_o({n7, n5}) );
endmodule


module flipflop_BITS1_22 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_22 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_22 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter2_4 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [1:0] request;
  output [1:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   tail_en, n1, n2;
  wire   [1:0] req_i;
  wire   [1:0] req_o;

  AND3X1 U10 ( .IN1(request[1]), .IN2(n1), .IN3(n2), .Q(grant[1]) );
  AND3X1 U11 ( .IN1(request[0]), .IN2(n2), .IN3(request[1]), .Q(tail_en) );
  INVX0 U6 ( .INP(request[0]), .ZN(n1) );
  NOR2X0 U7 ( .IN1(buffer_full_i), .IN2(n1), .QN(grant[0]) );
  INVX0 U8 ( .INP(buffer_full_i), .ZN(n2) );
  OA21X1 U9 ( .IN1(request[1]), .IN2(request[0]), .IN3(n2), .Q(grant_v_o) );
  register_BITS2_4 req_record ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i({1'b1, 1'b0}), .data_o({1'b0, 1'b0}) );
  register_BITS1_22 tail ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i(1'b1), .data_o(1'b0) );
endmodule


module flipflop_BITS4_26 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_26 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_26 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS4_25 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_25 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_25 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS4_24 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_24 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_24 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS1_21 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_21 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_21 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_20 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_20 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_20 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter4_8 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [3:0] request;
  output [3:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[2][3] , \req_i[2][2] , \req_i[2][1] , \req_i[2][0] ,
         \req_i[1][3] , \req_i[1][2] , \req_i[1][1] , \req_i[1][0] ,
         \req_i[0][3] , \req_i[0][2] , \req_i[0][1] , tail_en, N71, N265, N266,
         N267, N268, N276, N282, N291, N300, N301, N302, N303, n1, n2, n3, n4,
         n6, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21;
  wire   [2:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N265 = request[0];
  assign N266 = request[1];
  assign N267 = request[2];
  assign N268 = request[3];

  LATCHX1 shift_reg ( .CLK(1'b0), .D(1'b0), .Q(N71) );
  LATCHX1 \grant_reg[3]  ( .CLK(1'b1), .D(N303), .Q(grant[3]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N302), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N301), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N300), .Q(grant[0]) );
  LNANDX1 \req_i_reg[2][3]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][3] ) );
  LNANDX1 \req_i_reg[2][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][2] ) );
  LNANDX1 \req_i_reg[2][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][1] ) );
  LNANDX1 \req_i_reg[2][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][0] ) );
  LNANDX1 \req_i_reg[1][3]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][3] ) );
  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][3]  ( .CLK(tail_en), .D(N282), .Q(\req_i[0][3] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(n1), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(n4), .Q(\req_i[0][1] ) );
  LATCHX1 \tail_i_reg[0]  ( .CLK(tail_en), .D(N276), .Q(tail_i[0]) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N291), .D(tail_en), .Q(req_en[0]) );
  AND3X1 U35 ( .IN1(grant_v_o), .IN2(n19), .IN3(N267), .Q(N302) );
  NAND4X0 U37 ( .IN1(n17), .IN2(grant_v_o), .IN3(n16), .IN4(n20), .QN(N291) );
  AO21X1 U38 ( .IN1(n14), .IN2(n19), .IN3(buffer_full_i), .Q(n21) );
  NOR3X0 U39 ( .IN1(n4), .IN2(N282), .IN3(n1), .QN(n17) );
  NAND4X0 U41 ( .IN1(n11), .IN2(n13), .IN3(n9), .IN4(n10), .QN(N276) );
  AOI22X1 U42 ( .IN1(n2), .IN2(n15), .IN3(n15), .IN4(N265), .QN(n13) );
  AND2X1 U43 ( .IN1(N268), .IN2(n6), .Q(n15) );
  OA22X1 U44 ( .IN1(n6), .IN2(n18), .IN3(n6), .IN4(n3), .Q(n11) );
  INVX0 U15 ( .INP(N267), .ZN(n6) );
  INVX0 U16 ( .INP(n18), .ZN(n2) );
  NAND2X1 U17 ( .IN1(N266), .IN2(N265), .QN(n10) );
  NAND2X1 U18 ( .IN1(N267), .IN2(N268), .QN(n12) );
  INVX0 U19 ( .INP(N265), .ZN(n3) );
  NAND2X1 U20 ( .IN1(N266), .IN2(n3), .QN(n18) );
  NOR2X0 U21 ( .IN1(N266), .IN2(N265), .QN(n19) );
  INVX0 U22 ( .INP(n21), .ZN(grant_v_o) );
  NOR2X0 U23 ( .IN1(N268), .IN2(N267), .QN(n14) );
  NAND2X1 U24 ( .IN1(n15), .IN2(n19), .QN(n20) );
  NOR2X0 U25 ( .IN1(N265), .IN2(n2), .QN(n16) );
  NAND2X1 U26 ( .IN1(N71), .IN2(n7), .QN(n9) );
  INVX0 U27 ( .INP(n12), .ZN(n7) );
  INVX0 U28 ( .INP(n10), .ZN(n4) );
  INVX0 U29 ( .INP(n11), .ZN(n1) );
  NAND2X1 U30 ( .IN1(n13), .IN2(n12), .QN(N282) );
  NOR2X0 U31 ( .IN1(n21), .IN2(n17), .QN(tail_en) );
  NOR2X0 U32 ( .IN1(n3), .IN2(n21), .QN(N300) );
  NOR2X0 U33 ( .IN1(n18), .IN2(n21), .QN(N301) );
  NOR2X0 U34 ( .IN1(n21), .IN2(n20), .QN(N303) );
  register_BITS4_26 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][3] , \req_i[0][2] , \req_i[0][1] , 
        1'b0}), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS4_25 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][3] , \req_i[1][2] , \req_i[1][1] , 
        \req_i[1][0] }), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS4_24 \genblk1[2].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[2][3] , \req_i[2][2] , \req_i[2][1] , 
        \req_i[2][0] }), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS1_21 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(tail_i[0]), .data_o(1'b0) );
  register_BITS1_20 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module flipflop_BITS4_23 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_23 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_23 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS4_22 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_22 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_22 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS4_21 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_21 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_21 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS1_19 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_19 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_19 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_18 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_18 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_18 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter4_7 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [3:0] request;
  output [3:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[2][3] , \req_i[2][2] , \req_i[2][1] , \req_i[2][0] ,
         \req_i[1][3] , \req_i[1][2] , \req_i[1][1] , \req_i[1][0] ,
         \req_i[0][3] , \req_i[0][2] , \req_i[0][1] , tail_en, N71, N265, N266,
         N267, N268, N276, N282, N291, N300, N301, N302, N303, n1, n2, n3, n4,
         n6, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21;
  wire   [2:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N265 = request[0];
  assign N266 = request[1];
  assign N267 = request[2];
  assign N268 = request[3];

  LATCHX1 shift_reg ( .CLK(1'b0), .D(1'b0), .Q(N71) );
  LATCHX1 \grant_reg[3]  ( .CLK(1'b1), .D(N303), .Q(grant[3]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N302), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N301), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N300), .Q(grant[0]) );
  LNANDX1 \req_i_reg[2][3]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][3] ) );
  LNANDX1 \req_i_reg[2][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][2] ) );
  LNANDX1 \req_i_reg[2][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][1] ) );
  LNANDX1 \req_i_reg[2][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][0] ) );
  LNANDX1 \req_i_reg[1][3]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][3] ) );
  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][3]  ( .CLK(tail_en), .D(N282), .Q(\req_i[0][3] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(n1), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(n4), .Q(\req_i[0][1] ) );
  LATCHX1 \tail_i_reg[0]  ( .CLK(tail_en), .D(N276), .Q(tail_i[0]) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N291), .D(tail_en), .Q(req_en[0]) );
  AND3X1 U35 ( .IN1(grant_v_o), .IN2(n19), .IN3(N267), .Q(N302) );
  NAND4X0 U37 ( .IN1(n17), .IN2(grant_v_o), .IN3(n16), .IN4(n20), .QN(N291) );
  AO21X1 U38 ( .IN1(n14), .IN2(n19), .IN3(buffer_full_i), .Q(n21) );
  NOR3X0 U39 ( .IN1(n4), .IN2(N282), .IN3(n1), .QN(n17) );
  NAND4X0 U41 ( .IN1(n11), .IN2(n13), .IN3(n9), .IN4(n10), .QN(N276) );
  AOI22X1 U42 ( .IN1(n2), .IN2(n15), .IN3(n15), .IN4(N265), .QN(n13) );
  AND2X1 U43 ( .IN1(N268), .IN2(n6), .Q(n15) );
  OA22X1 U44 ( .IN1(n6), .IN2(n18), .IN3(n6), .IN4(n3), .Q(n11) );
  INVX0 U15 ( .INP(N267), .ZN(n6) );
  INVX0 U16 ( .INP(n18), .ZN(n2) );
  NAND2X1 U17 ( .IN1(N266), .IN2(N265), .QN(n10) );
  NAND2X1 U18 ( .IN1(N267), .IN2(N268), .QN(n12) );
  INVX0 U19 ( .INP(N265), .ZN(n3) );
  NAND2X1 U20 ( .IN1(N266), .IN2(n3), .QN(n18) );
  NOR2X0 U21 ( .IN1(N266), .IN2(N265), .QN(n19) );
  INVX0 U22 ( .INP(n21), .ZN(grant_v_o) );
  NOR2X0 U23 ( .IN1(N268), .IN2(N267), .QN(n14) );
  NAND2X1 U24 ( .IN1(n15), .IN2(n19), .QN(n20) );
  NOR2X0 U25 ( .IN1(N265), .IN2(n2), .QN(n16) );
  NAND2X1 U26 ( .IN1(N71), .IN2(n7), .QN(n9) );
  INVX0 U27 ( .INP(n12), .ZN(n7) );
  INVX0 U28 ( .INP(n10), .ZN(n4) );
  INVX0 U29 ( .INP(n11), .ZN(n1) );
  NAND2X1 U30 ( .IN1(n13), .IN2(n12), .QN(N282) );
  NOR2X0 U31 ( .IN1(n21), .IN2(n17), .QN(tail_en) );
  NOR2X0 U32 ( .IN1(n3), .IN2(n21), .QN(N300) );
  NOR2X0 U33 ( .IN1(n18), .IN2(n21), .QN(N301) );
  NOR2X0 U34 ( .IN1(n21), .IN2(n20), .QN(N303) );
  register_BITS4_23 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][3] , \req_i[0][2] , \req_i[0][1] , 
        1'b0}), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS4_22 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][3] , \req_i[1][2] , \req_i[1][1] , 
        \req_i[1][0] }), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS4_21 \genblk1[2].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[2][3] , \req_i[2][2] , \req_i[2][1] , 
        \req_i[2][0] }), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS1_19 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(tail_i[0]), .data_o(1'b0) );
  register_BITS1_18 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module flipflop_BITS4_20 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_20 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_20 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS4_19 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_19 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_19 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS4_18 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_18 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_18 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS1_17 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_17 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_17 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_16 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_16 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_16 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter4_6 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [3:0] request;
  output [3:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[2][3] , \req_i[2][2] , \req_i[2][1] , \req_i[2][0] ,
         \req_i[1][3] , \req_i[1][2] , \req_i[1][1] , \req_i[1][0] ,
         \req_i[0][3] , \req_i[0][2] , \req_i[0][1] , tail_en, N71, N265, N266,
         N267, N268, N276, N282, N291, N300, N301, N302, N303, n1, n2, n3, n4,
         n6, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21;
  wire   [2:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N265 = request[0];
  assign N266 = request[1];
  assign N267 = request[2];
  assign N268 = request[3];

  LATCHX1 shift_reg ( .CLK(1'b0), .D(1'b0), .Q(N71) );
  LATCHX1 \grant_reg[3]  ( .CLK(1'b1), .D(N303), .Q(grant[3]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N302), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N301), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N300), .Q(grant[0]) );
  LNANDX1 \req_i_reg[2][3]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][3] ) );
  LNANDX1 \req_i_reg[2][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][2] ) );
  LNANDX1 \req_i_reg[2][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][1] ) );
  LNANDX1 \req_i_reg[2][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][0] ) );
  LNANDX1 \req_i_reg[1][3]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][3] ) );
  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][3]  ( .CLK(tail_en), .D(N282), .Q(\req_i[0][3] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(n1), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(n4), .Q(\req_i[0][1] ) );
  LATCHX1 \tail_i_reg[0]  ( .CLK(tail_en), .D(N276), .Q(tail_i[0]) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N291), .D(tail_en), .Q(req_en[0]) );
  AND3X1 U35 ( .IN1(grant_v_o), .IN2(n19), .IN3(N267), .Q(N302) );
  NAND4X0 U37 ( .IN1(n17), .IN2(grant_v_o), .IN3(n16), .IN4(n20), .QN(N291) );
  AO21X1 U38 ( .IN1(n14), .IN2(n19), .IN3(buffer_full_i), .Q(n21) );
  NOR3X0 U39 ( .IN1(n4), .IN2(N282), .IN3(n1), .QN(n17) );
  NAND4X0 U41 ( .IN1(n11), .IN2(n13), .IN3(n9), .IN4(n10), .QN(N276) );
  AOI22X1 U42 ( .IN1(n2), .IN2(n15), .IN3(n15), .IN4(N265), .QN(n13) );
  AND2X1 U43 ( .IN1(N268), .IN2(n6), .Q(n15) );
  OA22X1 U44 ( .IN1(n6), .IN2(n18), .IN3(n6), .IN4(n3), .Q(n11) );
  INVX0 U15 ( .INP(N267), .ZN(n6) );
  INVX0 U16 ( .INP(n18), .ZN(n2) );
  NAND2X1 U17 ( .IN1(N266), .IN2(N265), .QN(n10) );
  NAND2X1 U18 ( .IN1(N267), .IN2(N268), .QN(n12) );
  INVX0 U19 ( .INP(N265), .ZN(n3) );
  NAND2X1 U20 ( .IN1(N266), .IN2(n3), .QN(n18) );
  NOR2X0 U21 ( .IN1(N266), .IN2(N265), .QN(n19) );
  INVX0 U22 ( .INP(n21), .ZN(grant_v_o) );
  NOR2X0 U23 ( .IN1(N268), .IN2(N267), .QN(n14) );
  NAND2X1 U24 ( .IN1(n15), .IN2(n19), .QN(n20) );
  NOR2X0 U25 ( .IN1(N265), .IN2(n2), .QN(n16) );
  NAND2X1 U26 ( .IN1(N71), .IN2(n7), .QN(n9) );
  INVX0 U27 ( .INP(n12), .ZN(n7) );
  INVX0 U28 ( .INP(n10), .ZN(n4) );
  INVX0 U29 ( .INP(n11), .ZN(n1) );
  NAND2X1 U30 ( .IN1(n13), .IN2(n12), .QN(N282) );
  NOR2X0 U31 ( .IN1(n21), .IN2(n17), .QN(tail_en) );
  NOR2X0 U32 ( .IN1(n3), .IN2(n21), .QN(N300) );
  NOR2X0 U33 ( .IN1(n18), .IN2(n21), .QN(N301) );
  NOR2X0 U34 ( .IN1(n21), .IN2(n20), .QN(N303) );
  register_BITS4_20 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][3] , \req_i[0][2] , \req_i[0][1] , 
        1'b0}), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS4_19 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][3] , \req_i[1][2] , \req_i[1][1] , 
        \req_i[1][0] }), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS4_18 \genblk1[2].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[2][3] , \req_i[2][2] , \req_i[2][1] , 
        \req_i[2][0] }), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS1_17 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(tail_i[0]), .data_o(1'b0) );
  register_BITS1_16 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module dccl_14 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_13 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_12 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_11 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_10 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module controller5_2 ( clk, rst, .packet_addr({\packet_addr[4][7] , 
        \packet_addr[4][6] , \packet_addr[4][5] , \packet_addr[4][4] , 
        \packet_addr[4][3] , \packet_addr[4][2] , \packet_addr[4][1] , 
        \packet_addr[4][0] , \packet_addr[3][7] , \packet_addr[3][6] , 
        \packet_addr[3][5] , \packet_addr[3][4] , \packet_addr[3][3] , 
        \packet_addr[3][2] , \packet_addr[3][1] , \packet_addr[3][0] , 
        \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] , 
        \packet_addr[2][4] , \packet_addr[2][3] , \packet_addr[2][2] , 
        \packet_addr[2][1] , \packet_addr[2][0] , \packet_addr[1][7] , 
        \packet_addr[1][6] , \packet_addr[1][5] , \packet_addr[1][4] , 
        \packet_addr[1][3] , \packet_addr[1][2] , \packet_addr[1][1] , 
        \packet_addr[1][0] , \packet_addr[0][7] , \packet_addr[0][6] , 
        \packet_addr[0][5] , \packet_addr[0][4] , \packet_addr[0][3] , 
        \packet_addr[0][2] , \packet_addr[0][1] , \packet_addr[0][0] }), 
        local_addr, packet_valid, buffer_full_in, grant_0, grant_1, grant_2, 
        grant_3, grant_4, grant_v, pop_v );
  input [7:0] local_addr;
  input [4:0] packet_valid;
  input [4:0] buffer_full_in;
  output [1:0] grant_0;
  output [1:0] grant_1;
  output [3:0] grant_2;
  output [3:0] grant_3;
  output [3:0] grant_4;
  output [4:0] grant_v;
  output [4:0] pop_v;
  input clk, rst, \packet_addr[4][7] , \packet_addr[4][6] ,
         \packet_addr[4][5] , \packet_addr[4][4] , \packet_addr[4][3] ,
         \packet_addr[4][2] , \packet_addr[4][1] , \packet_addr[4][0] ,
         \packet_addr[3][7] , \packet_addr[3][6] , \packet_addr[3][5] ,
         \packet_addr[3][4] , \packet_addr[3][3] , \packet_addr[3][2] ,
         \packet_addr[3][1] , \packet_addr[3][0] , \packet_addr[2][7] ,
         \packet_addr[2][6] , \packet_addr[2][5] , \packet_addr[2][4] ,
         \packet_addr[2][3] , \packet_addr[2][2] , \packet_addr[2][1] ,
         \packet_addr[2][0] , \packet_addr[1][7] , \packet_addr[1][6] ,
         \packet_addr[1][5] , \packet_addr[1][4] , \packet_addr[1][3] ,
         \packet_addr[1][2] , \packet_addr[1][1] , \packet_addr[1][0] ,
         \packet_addr[0][7] , \packet_addr[0][6] , \packet_addr[0][5] ,
         \packet_addr[0][4] , \packet_addr[0][3] , \packet_addr[0][2] ,
         \packet_addr[0][1] , \packet_addr[0][0] ;
  wire   \request[4][3] , \request[4][2] , \request[4][1] , \request[4][0] ,
         \request[3][3] , \request[3][2] , \request[3][1] , \request[3][0] ,
         \request[2][3] , \request[2][2] , \request[2][1] , \request[2][0] ,
         \request[1][1] , \request[1][0] , \request[0][1] , \request[0][0] ;

  OR4X1 U1 ( .IN1(grant_1[1]), .IN2(grant_0[1]), .IN3(grant_3[3]), .IN4(
        grant_2[3]), .Q(pop_v[4]) );
  OR2X1 U2 ( .IN1(grant_2[2]), .IN2(grant_4[3]), .Q(pop_v[3]) );
  OR2X1 U3 ( .IN1(grant_3[2]), .IN2(grant_4[2]), .Q(pop_v[2]) );
  OR4X1 U4 ( .IN1(grant_2[1]), .IN2(grant_0[0]), .IN3(grant_4[1]), .IN4(
        grant_3[1]), .Q(pop_v[1]) );
  OR4X1 U5 ( .IN1(grant_2[0]), .IN2(grant_1[0]), .IN3(grant_4[0]), .IN4(
        grant_3[0]), .Q(pop_v[0]) );
  arbiter2_5 arbiter_n ( .clk(clk), .rst(rst), .request({\request[0][1] , 
        \request[0][0] }), .buffer_full_i(buffer_full_in[0]), .grant(grant_0), 
        .grant_v_o(grant_v[0]) );
  arbiter2_4 arbiter_s ( .clk(clk), .rst(rst), .request({\request[1][1] , 
        \request[1][0] }), .buffer_full_i(buffer_full_in[1]), .grant(grant_1), 
        .grant_v_o(grant_v[1]) );
  arbiter4_8 arbiter_e ( .clk(clk), .rst(rst), .request({\request[2][3] , 
        \request[2][2] , \request[2][1] , \request[2][0] }), .buffer_full_i(
        buffer_full_in[2]), .grant(grant_2), .grant_v_o(grant_v[2]) );
  arbiter4_7 arbiter_w ( .clk(clk), .rst(rst), .request({\request[3][3] , 
        \request[3][2] , \request[3][1] , \request[3][0] }), .buffer_full_i(
        buffer_full_in[3]), .grant(grant_3), .grant_v_o(grant_v[3]) );
  arbiter4_6 arbiter_l ( .clk(clk), .rst(rst), .request({\request[4][3] , 
        \request[4][2] , \request[4][1] , \request[4][0] }), .buffer_full_i(
        buffer_full_in[4]), .grant(grant_4), .grant_v_o(grant_v[4]) );
  dccl_14 dccl_n ( .packet_addr_y_i({\packet_addr[0][3] , \packet_addr[0][2] , 
        \packet_addr[0][1] , \packet_addr[0][0] }), .packet_addr_x_i({
        \packet_addr[0][7] , \packet_addr[0][6] , \packet_addr[0][5] , 
        \packet_addr[0][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[0]), 
        .east_req(\request[2][0] ), .south_req(\request[1][0] ), .west_req(
        \request[3][0] ), .local_req(\request[4][0] ) );
  dccl_13 dccl_s ( .packet_addr_y_i({\packet_addr[1][3] , \packet_addr[1][2] , 
        \packet_addr[1][1] , \packet_addr[1][0] }), .packet_addr_x_i({
        \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] , 
        \packet_addr[1][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[1]), 
        .north_req(\request[0][0] ), .east_req(\request[2][1] ), .west_req(
        \request[3][1] ), .local_req(\request[4][1] ) );
  dccl_12 dccl_e ( .packet_addr_y_i({\packet_addr[2][3] , \packet_addr[2][2] , 
        \packet_addr[2][1] , \packet_addr[2][0] }), .packet_addr_x_i({
        \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] , 
        \packet_addr[2][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[2]), 
        .west_req(\request[3][2] ), .local_req(\request[4][2] ) );
  dccl_11 dccl_w ( .packet_addr_y_i({\packet_addr[3][3] , \packet_addr[3][2] , 
        \packet_addr[3][1] , \packet_addr[3][0] }), .packet_addr_x_i({
        \packet_addr[3][7] , \packet_addr[3][6] , \packet_addr[3][5] , 
        \packet_addr[3][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[3]), 
        .east_req(\request[2][2] ), .local_req(\request[4][3] ) );
  dccl_10 dccl_l ( .packet_addr_y_i({\packet_addr[4][3] , \packet_addr[4][2] , 
        \packet_addr[4][1] , \packet_addr[4][0] }), .packet_addr_x_i({
        \packet_addr[4][7] , \packet_addr[4][6] , \packet_addr[4][5] , 
        \packet_addr[4][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[4]), 
        .north_req(\request[0][1] ), .east_req(\request[2][3] ), .south_req(
        \request[1][1] ), .west_req(\request[3][3] ) );
endmodule


module mux2_1_5 ( data0, data1, select0, select1, data_o );
  input [15:0] data0;
  input [15:0] data1;
  output [15:0] data_o;
  input select0, select1;
  wire   n1, n4, n5;

  AO22X1 U4 ( .IN1(data1[9]), .IN2(n5), .IN3(data0[9]), .IN4(n4), .Q(data_o[9]) );
  AO22X1 U5 ( .IN1(data1[8]), .IN2(n5), .IN3(data0[8]), .IN4(n4), .Q(data_o[8]) );
  AO22X1 U6 ( .IN1(data1[7]), .IN2(n5), .IN3(data0[7]), .IN4(n4), .Q(data_o[7]) );
  AO22X1 U7 ( .IN1(data1[6]), .IN2(n5), .IN3(data0[6]), .IN4(n4), .Q(data_o[6]) );
  AO22X1 U8 ( .IN1(data1[5]), .IN2(n5), .IN3(data0[5]), .IN4(n4), .Q(data_o[5]) );
  AO22X1 U9 ( .IN1(data1[4]), .IN2(n5), .IN3(data0[4]), .IN4(n4), .Q(data_o[4]) );
  AO22X1 U10 ( .IN1(data1[3]), .IN2(n5), .IN3(data0[3]), .IN4(n4), .Q(
        data_o[3]) );
  AO22X1 U11 ( .IN1(data1[2]), .IN2(n5), .IN3(data0[2]), .IN4(n4), .Q(
        data_o[2]) );
  AO22X1 U12 ( .IN1(data1[1]), .IN2(n5), .IN3(data0[1]), .IN4(n4), .Q(
        data_o[1]) );
  AO22X1 U13 ( .IN1(data1[15]), .IN2(n5), .IN3(data0[15]), .IN4(n4), .Q(
        data_o[15]) );
  AO22X1 U14 ( .IN1(data1[14]), .IN2(n5), .IN3(data0[14]), .IN4(n4), .Q(
        data_o[14]) );
  AO22X1 U15 ( .IN1(data1[13]), .IN2(n5), .IN3(data0[13]), .IN4(n4), .Q(
        data_o[13]) );
  AO22X1 U16 ( .IN1(data1[12]), .IN2(n5), .IN3(data0[12]), .IN4(n4), .Q(
        data_o[12]) );
  AO22X1 U17 ( .IN1(data1[11]), .IN2(n5), .IN3(data0[11]), .IN4(n4), .Q(
        data_o[11]) );
  AO22X1 U18 ( .IN1(data1[10]), .IN2(n5), .IN3(data0[10]), .IN4(n4), .Q(
        data_o[10]) );
  AO22X1 U19 ( .IN1(data1[0]), .IN2(n5), .IN3(data0[0]), .IN4(n4), .Q(
        data_o[0]) );
  INVX0 U2 ( .INP(select1), .ZN(n1) );
  AND2X1 U3 ( .IN1(select0), .IN2(n1), .Q(n4) );
  NOR2X0 U20 ( .IN1(n1), .IN2(select0), .QN(n5) );
endmodule


module mux2_1_4 ( data0, data1, select0, select1, data_o );
  input [15:0] data0;
  input [15:0] data1;
  output [15:0] data_o;
  input select0, select1;
  wire   n1, n4, n5;

  AO22X1 U4 ( .IN1(data1[9]), .IN2(n5), .IN3(data0[9]), .IN4(n4), .Q(data_o[9]) );
  AO22X1 U5 ( .IN1(data1[8]), .IN2(n5), .IN3(data0[8]), .IN4(n4), .Q(data_o[8]) );
  AO22X1 U6 ( .IN1(data1[7]), .IN2(n5), .IN3(data0[7]), .IN4(n4), .Q(data_o[7]) );
  AO22X1 U7 ( .IN1(data1[6]), .IN2(n5), .IN3(data0[6]), .IN4(n4), .Q(data_o[6]) );
  AO22X1 U8 ( .IN1(data1[5]), .IN2(n5), .IN3(data0[5]), .IN4(n4), .Q(data_o[5]) );
  AO22X1 U9 ( .IN1(data1[4]), .IN2(n5), .IN3(data0[4]), .IN4(n4), .Q(data_o[4]) );
  AO22X1 U10 ( .IN1(data1[3]), .IN2(n5), .IN3(data0[3]), .IN4(n4), .Q(
        data_o[3]) );
  AO22X1 U11 ( .IN1(data1[2]), .IN2(n5), .IN3(data0[2]), .IN4(n4), .Q(
        data_o[2]) );
  AO22X1 U12 ( .IN1(data1[1]), .IN2(n5), .IN3(data0[1]), .IN4(n4), .Q(
        data_o[1]) );
  AO22X1 U13 ( .IN1(data1[15]), .IN2(n5), .IN3(data0[15]), .IN4(n4), .Q(
        data_o[15]) );
  AO22X1 U14 ( .IN1(data1[14]), .IN2(n5), .IN3(data0[14]), .IN4(n4), .Q(
        data_o[14]) );
  AO22X1 U15 ( .IN1(data1[13]), .IN2(n5), .IN3(data0[13]), .IN4(n4), .Q(
        data_o[13]) );
  AO22X1 U16 ( .IN1(data1[12]), .IN2(n5), .IN3(data0[12]), .IN4(n4), .Q(
        data_o[12]) );
  AO22X1 U17 ( .IN1(data1[11]), .IN2(n5), .IN3(data0[11]), .IN4(n4), .Q(
        data_o[11]) );
  AO22X1 U18 ( .IN1(data1[10]), .IN2(n5), .IN3(data0[10]), .IN4(n4), .Q(
        data_o[10]) );
  AO22X1 U19 ( .IN1(data1[0]), .IN2(n5), .IN3(data0[0]), .IN4(n4), .Q(
        data_o[0]) );
  INVX0 U2 ( .INP(select1), .ZN(n1) );
  AND2X1 U3 ( .IN1(select0), .IN2(n1), .Q(n4) );
  NOR2X0 U20 ( .IN1(n1), .IN2(select0), .QN(n5) );
endmodule


module mux4_1_8 ( data0, data1, data2, data3, select0, select1, select2, 
        select3, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  input [15:0] data3;
  output [15:0] data_o;
  input select0, select1, select2, select3;
  wire   n1, n2, n3, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43;

  AO221X1 U5 ( .IN1(data1[9]), .IN2(n43), .IN3(data0[9]), .IN4(n42), .IN5(n41), 
        .Q(data_o[9]) );
  AO22X1 U6 ( .IN1(data2[9]), .IN2(n40), .IN3(data3[9]), .IN4(n39), .Q(n41) );
  AO221X1 U7 ( .IN1(data1[8]), .IN2(n43), .IN3(data0[8]), .IN4(n42), .IN5(n38), 
        .Q(data_o[8]) );
  AO22X1 U8 ( .IN1(data2[8]), .IN2(n40), .IN3(data3[8]), .IN4(n39), .Q(n38) );
  AO221X1 U9 ( .IN1(data1[7]), .IN2(n43), .IN3(data0[7]), .IN4(n42), .IN5(n37), 
        .Q(data_o[7]) );
  AO22X1 U10 ( .IN1(data2[7]), .IN2(n40), .IN3(data3[7]), .IN4(n39), .Q(n37)
         );
  AO221X1 U11 ( .IN1(data1[6]), .IN2(n43), .IN3(data0[6]), .IN4(n42), .IN5(n36), .Q(data_o[6]) );
  AO22X1 U12 ( .IN1(data2[6]), .IN2(n40), .IN3(data3[6]), .IN4(n39), .Q(n36)
         );
  AO221X1 U13 ( .IN1(data1[5]), .IN2(n43), .IN3(data0[5]), .IN4(n42), .IN5(n35), .Q(data_o[5]) );
  AO22X1 U14 ( .IN1(data2[5]), .IN2(n40), .IN3(data3[5]), .IN4(n39), .Q(n35)
         );
  AO221X1 U15 ( .IN1(data1[4]), .IN2(n43), .IN3(data0[4]), .IN4(n42), .IN5(n34), .Q(data_o[4]) );
  AO22X1 U16 ( .IN1(data2[4]), .IN2(n40), .IN3(data3[4]), .IN4(n39), .Q(n34)
         );
  AO221X1 U17 ( .IN1(data1[3]), .IN2(n43), .IN3(data0[3]), .IN4(n42), .IN5(n33), .Q(data_o[3]) );
  AO22X1 U18 ( .IN1(data2[3]), .IN2(n40), .IN3(data3[3]), .IN4(n39), .Q(n33)
         );
  AO221X1 U19 ( .IN1(data1[2]), .IN2(n43), .IN3(data0[2]), .IN4(n42), .IN5(n32), .Q(data_o[2]) );
  AO22X1 U20 ( .IN1(data2[2]), .IN2(n40), .IN3(data3[2]), .IN4(n39), .Q(n32)
         );
  AO221X1 U21 ( .IN1(data1[1]), .IN2(n43), .IN3(data0[1]), .IN4(n42), .IN5(n31), .Q(data_o[1]) );
  AO22X1 U22 ( .IN1(data2[1]), .IN2(n40), .IN3(data3[1]), .IN4(n39), .Q(n31)
         );
  AO221X1 U23 ( .IN1(data1[15]), .IN2(n43), .IN3(data0[15]), .IN4(n42), .IN5(
        n30), .Q(data_o[15]) );
  AO22X1 U24 ( .IN1(data2[15]), .IN2(n40), .IN3(data3[15]), .IN4(n39), .Q(n30)
         );
  AO221X1 U25 ( .IN1(data1[14]), .IN2(n43), .IN3(data0[14]), .IN4(n42), .IN5(
        n29), .Q(data_o[14]) );
  AO22X1 U26 ( .IN1(data2[14]), .IN2(n40), .IN3(data3[14]), .IN4(n39), .Q(n29)
         );
  AO221X1 U27 ( .IN1(data1[13]), .IN2(n43), .IN3(data0[13]), .IN4(n42), .IN5(
        n28), .Q(data_o[13]) );
  AO22X1 U28 ( .IN1(data2[13]), .IN2(n40), .IN3(data3[13]), .IN4(n39), .Q(n28)
         );
  AO221X1 U29 ( .IN1(data1[12]), .IN2(n43), .IN3(data0[12]), .IN4(n42), .IN5(
        n27), .Q(data_o[12]) );
  AO22X1 U30 ( .IN1(data2[12]), .IN2(n40), .IN3(data3[12]), .IN4(n39), .Q(n27)
         );
  AO221X1 U31 ( .IN1(data1[11]), .IN2(n43), .IN3(data0[11]), .IN4(n42), .IN5(
        n26), .Q(data_o[11]) );
  AO22X1 U32 ( .IN1(data2[11]), .IN2(n40), .IN3(data3[11]), .IN4(n39), .Q(n26)
         );
  AO221X1 U33 ( .IN1(data1[10]), .IN2(n43), .IN3(data0[10]), .IN4(n42), .IN5(
        n25), .Q(data_o[10]) );
  AO22X1 U34 ( .IN1(data2[10]), .IN2(n40), .IN3(data3[10]), .IN4(n39), .Q(n25)
         );
  AO221X1 U35 ( .IN1(data1[0]), .IN2(n43), .IN3(data0[0]), .IN4(n42), .IN5(n24), .Q(data_o[0]) );
  AO22X1 U36 ( .IN1(data2[0]), .IN2(n40), .IN3(data3[0]), .IN4(n39), .Q(n24)
         );
  INVX0 U2 ( .INP(select2), .ZN(n1) );
  NOR4X0 U3 ( .IN1(n1), .IN2(select0), .IN3(select1), .IN4(select3), .QN(n40)
         );
  AND4X1 U4 ( .IN1(select3), .IN2(n3), .IN3(n2), .IN4(n1), .Q(n39) );
  INVX0 U37 ( .INP(select0), .ZN(n3) );
  INVX0 U38 ( .INP(select1), .ZN(n2) );
  NOR4X0 U39 ( .IN1(n3), .IN2(select1), .IN3(select2), .IN4(select3), .QN(n42)
         );
  NOR4X0 U40 ( .IN1(n2), .IN2(select0), .IN3(select2), .IN4(select3), .QN(n43)
         );
endmodule


module mux4_1_7 ( data0, data1, data2, data3, select0, select1, select2, 
        select3, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  input [15:0] data3;
  output [15:0] data_o;
  input select0, select1, select2, select3;
  wire   n1, n2, n3, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43;

  AO221X1 U5 ( .IN1(data1[9]), .IN2(n43), .IN3(data0[9]), .IN4(n42), .IN5(n41), 
        .Q(data_o[9]) );
  AO22X1 U6 ( .IN1(data2[9]), .IN2(n40), .IN3(data3[9]), .IN4(n39), .Q(n41) );
  AO221X1 U7 ( .IN1(data1[8]), .IN2(n43), .IN3(data0[8]), .IN4(n42), .IN5(n38), 
        .Q(data_o[8]) );
  AO22X1 U8 ( .IN1(data2[8]), .IN2(n40), .IN3(data3[8]), .IN4(n39), .Q(n38) );
  AO221X1 U9 ( .IN1(data1[7]), .IN2(n43), .IN3(data0[7]), .IN4(n42), .IN5(n37), 
        .Q(data_o[7]) );
  AO22X1 U10 ( .IN1(data2[7]), .IN2(n40), .IN3(data3[7]), .IN4(n39), .Q(n37)
         );
  AO221X1 U11 ( .IN1(data1[6]), .IN2(n43), .IN3(data0[6]), .IN4(n42), .IN5(n36), .Q(data_o[6]) );
  AO22X1 U12 ( .IN1(data2[6]), .IN2(n40), .IN3(data3[6]), .IN4(n39), .Q(n36)
         );
  AO221X1 U13 ( .IN1(data1[5]), .IN2(n43), .IN3(data0[5]), .IN4(n42), .IN5(n35), .Q(data_o[5]) );
  AO22X1 U14 ( .IN1(data2[5]), .IN2(n40), .IN3(data3[5]), .IN4(n39), .Q(n35)
         );
  AO221X1 U15 ( .IN1(data1[4]), .IN2(n43), .IN3(data0[4]), .IN4(n42), .IN5(n34), .Q(data_o[4]) );
  AO22X1 U16 ( .IN1(data2[4]), .IN2(n40), .IN3(data3[4]), .IN4(n39), .Q(n34)
         );
  AO221X1 U17 ( .IN1(data1[3]), .IN2(n43), .IN3(data0[3]), .IN4(n42), .IN5(n33), .Q(data_o[3]) );
  AO22X1 U18 ( .IN1(data2[3]), .IN2(n40), .IN3(data3[3]), .IN4(n39), .Q(n33)
         );
  AO221X1 U19 ( .IN1(data1[2]), .IN2(n43), .IN3(data0[2]), .IN4(n42), .IN5(n32), .Q(data_o[2]) );
  AO22X1 U20 ( .IN1(data2[2]), .IN2(n40), .IN3(data3[2]), .IN4(n39), .Q(n32)
         );
  AO221X1 U21 ( .IN1(data1[1]), .IN2(n43), .IN3(data0[1]), .IN4(n42), .IN5(n31), .Q(data_o[1]) );
  AO22X1 U22 ( .IN1(data2[1]), .IN2(n40), .IN3(data3[1]), .IN4(n39), .Q(n31)
         );
  AO221X1 U23 ( .IN1(data1[15]), .IN2(n43), .IN3(data0[15]), .IN4(n42), .IN5(
        n30), .Q(data_o[15]) );
  AO22X1 U24 ( .IN1(data2[15]), .IN2(n40), .IN3(data3[15]), .IN4(n39), .Q(n30)
         );
  AO221X1 U25 ( .IN1(data1[14]), .IN2(n43), .IN3(data0[14]), .IN4(n42), .IN5(
        n29), .Q(data_o[14]) );
  AO22X1 U26 ( .IN1(data2[14]), .IN2(n40), .IN3(data3[14]), .IN4(n39), .Q(n29)
         );
  AO221X1 U27 ( .IN1(data1[13]), .IN2(n43), .IN3(data0[13]), .IN4(n42), .IN5(
        n28), .Q(data_o[13]) );
  AO22X1 U28 ( .IN1(data2[13]), .IN2(n40), .IN3(data3[13]), .IN4(n39), .Q(n28)
         );
  AO221X1 U29 ( .IN1(data1[12]), .IN2(n43), .IN3(data0[12]), .IN4(n42), .IN5(
        n27), .Q(data_o[12]) );
  AO22X1 U30 ( .IN1(data2[12]), .IN2(n40), .IN3(data3[12]), .IN4(n39), .Q(n27)
         );
  AO221X1 U31 ( .IN1(data1[11]), .IN2(n43), .IN3(data0[11]), .IN4(n42), .IN5(
        n26), .Q(data_o[11]) );
  AO22X1 U32 ( .IN1(data2[11]), .IN2(n40), .IN3(data3[11]), .IN4(n39), .Q(n26)
         );
  AO221X1 U33 ( .IN1(data1[10]), .IN2(n43), .IN3(data0[10]), .IN4(n42), .IN5(
        n25), .Q(data_o[10]) );
  AO22X1 U34 ( .IN1(data2[10]), .IN2(n40), .IN3(data3[10]), .IN4(n39), .Q(n25)
         );
  AO221X1 U35 ( .IN1(data1[0]), .IN2(n43), .IN3(data0[0]), .IN4(n42), .IN5(n24), .Q(data_o[0]) );
  AO22X1 U36 ( .IN1(data2[0]), .IN2(n40), .IN3(data3[0]), .IN4(n39), .Q(n24)
         );
  INVX0 U2 ( .INP(select2), .ZN(n1) );
  NOR4X0 U3 ( .IN1(n1), .IN2(select0), .IN3(select1), .IN4(select3), .QN(n40)
         );
  AND4X1 U4 ( .IN1(select3), .IN2(n3), .IN3(n2), .IN4(n1), .Q(n39) );
  INVX0 U37 ( .INP(select0), .ZN(n3) );
  INVX0 U38 ( .INP(select1), .ZN(n2) );
  NOR4X0 U39 ( .IN1(n3), .IN2(select1), .IN3(select2), .IN4(select3), .QN(n42)
         );
  NOR4X0 U40 ( .IN1(n2), .IN2(select0), .IN3(select2), .IN4(select3), .QN(n43)
         );
endmodule


module mux4_1_6 ( data0, data1, data2, data3, select0, select1, select2, 
        select3, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  input [15:0] data3;
  output [15:0] data_o;
  input select0, select1, select2, select3;
  wire   n1, n2, n3, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43;

  AO221X1 U5 ( .IN1(data1[9]), .IN2(n43), .IN3(data0[9]), .IN4(n42), .IN5(n41), 
        .Q(data_o[9]) );
  AO22X1 U6 ( .IN1(data2[9]), .IN2(n40), .IN3(data3[9]), .IN4(n39), .Q(n41) );
  AO221X1 U7 ( .IN1(data1[8]), .IN2(n43), .IN3(data0[8]), .IN4(n42), .IN5(n38), 
        .Q(data_o[8]) );
  AO22X1 U8 ( .IN1(data2[8]), .IN2(n40), .IN3(data3[8]), .IN4(n39), .Q(n38) );
  AO221X1 U9 ( .IN1(data1[7]), .IN2(n43), .IN3(data0[7]), .IN4(n42), .IN5(n37), 
        .Q(data_o[7]) );
  AO22X1 U10 ( .IN1(data2[7]), .IN2(n40), .IN3(data3[7]), .IN4(n39), .Q(n37)
         );
  AO221X1 U11 ( .IN1(data1[6]), .IN2(n43), .IN3(data0[6]), .IN4(n42), .IN5(n36), .Q(data_o[6]) );
  AO22X1 U12 ( .IN1(data2[6]), .IN2(n40), .IN3(data3[6]), .IN4(n39), .Q(n36)
         );
  AO221X1 U13 ( .IN1(data1[5]), .IN2(n43), .IN3(data0[5]), .IN4(n42), .IN5(n35), .Q(data_o[5]) );
  AO22X1 U14 ( .IN1(data2[5]), .IN2(n40), .IN3(data3[5]), .IN4(n39), .Q(n35)
         );
  AO221X1 U15 ( .IN1(data1[4]), .IN2(n43), .IN3(data0[4]), .IN4(n42), .IN5(n34), .Q(data_o[4]) );
  AO22X1 U16 ( .IN1(data2[4]), .IN2(n40), .IN3(data3[4]), .IN4(n39), .Q(n34)
         );
  AO221X1 U17 ( .IN1(data1[3]), .IN2(n43), .IN3(data0[3]), .IN4(n42), .IN5(n33), .Q(data_o[3]) );
  AO22X1 U18 ( .IN1(data2[3]), .IN2(n40), .IN3(data3[3]), .IN4(n39), .Q(n33)
         );
  AO221X1 U19 ( .IN1(data1[2]), .IN2(n43), .IN3(data0[2]), .IN4(n42), .IN5(n32), .Q(data_o[2]) );
  AO22X1 U20 ( .IN1(data2[2]), .IN2(n40), .IN3(data3[2]), .IN4(n39), .Q(n32)
         );
  AO221X1 U21 ( .IN1(data1[1]), .IN2(n43), .IN3(data0[1]), .IN4(n42), .IN5(n31), .Q(data_o[1]) );
  AO22X1 U22 ( .IN1(data2[1]), .IN2(n40), .IN3(data3[1]), .IN4(n39), .Q(n31)
         );
  AO221X1 U23 ( .IN1(data1[15]), .IN2(n43), .IN3(data0[15]), .IN4(n42), .IN5(
        n30), .Q(data_o[15]) );
  AO22X1 U24 ( .IN1(data2[15]), .IN2(n40), .IN3(data3[15]), .IN4(n39), .Q(n30)
         );
  AO221X1 U25 ( .IN1(data1[14]), .IN2(n43), .IN3(data0[14]), .IN4(n42), .IN5(
        n29), .Q(data_o[14]) );
  AO22X1 U26 ( .IN1(data2[14]), .IN2(n40), .IN3(data3[14]), .IN4(n39), .Q(n29)
         );
  AO221X1 U27 ( .IN1(data1[13]), .IN2(n43), .IN3(data0[13]), .IN4(n42), .IN5(
        n28), .Q(data_o[13]) );
  AO22X1 U28 ( .IN1(data2[13]), .IN2(n40), .IN3(data3[13]), .IN4(n39), .Q(n28)
         );
  AO221X1 U29 ( .IN1(data1[12]), .IN2(n43), .IN3(data0[12]), .IN4(n42), .IN5(
        n27), .Q(data_o[12]) );
  AO22X1 U30 ( .IN1(data2[12]), .IN2(n40), .IN3(data3[12]), .IN4(n39), .Q(n27)
         );
  AO221X1 U31 ( .IN1(data1[11]), .IN2(n43), .IN3(data0[11]), .IN4(n42), .IN5(
        n26), .Q(data_o[11]) );
  AO22X1 U32 ( .IN1(data2[11]), .IN2(n40), .IN3(data3[11]), .IN4(n39), .Q(n26)
         );
  AO221X1 U33 ( .IN1(data1[10]), .IN2(n43), .IN3(data0[10]), .IN4(n42), .IN5(
        n25), .Q(data_o[10]) );
  AO22X1 U34 ( .IN1(data2[10]), .IN2(n40), .IN3(data3[10]), .IN4(n39), .Q(n25)
         );
  AO221X1 U35 ( .IN1(data1[0]), .IN2(n43), .IN3(data0[0]), .IN4(n42), .IN5(n24), .Q(data_o[0]) );
  AO22X1 U36 ( .IN1(data2[0]), .IN2(n40), .IN3(data3[0]), .IN4(n39), .Q(n24)
         );
  INVX0 U2 ( .INP(select2), .ZN(n1) );
  NOR4X0 U3 ( .IN1(n1), .IN2(select0), .IN3(select1), .IN4(select3), .QN(n40)
         );
  AND4X1 U4 ( .IN1(select3), .IN2(n3), .IN3(n2), .IN4(n1), .Q(n39) );
  INVX0 U37 ( .INP(select0), .ZN(n3) );
  INVX0 U38 ( .INP(select1), .ZN(n2) );
  NOR4X0 U39 ( .IN1(n3), .IN2(select1), .IN3(select2), .IN4(select3), .QN(n42)
         );
  NOR4X0 U40 ( .IN1(n2), .IN2(select0), .IN3(select2), .IN4(select3), .QN(n43)
         );
endmodule



    module node5_NODE_X1_NODE_Y2I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__I_node_2_node_interface__I_node_3_node_interface__ ( 
        \clk.clk , \reset.reset , \local_node.clk , 
        \local_node.buffer_full_in , \local_node.buffer_full_out , 
        \local_node.receiving_data , \local_node.sending_data , 
        \local_node.data_in , \local_node.data_out , \node_0.clk , 
        \node_0.buffer_full_in , \node_0.buffer_full_out , 
        \node_0.receiving_data , \node_0.sending_data , \node_0.data_in , 
        \node_0.data_out , \node_1.clk , \node_1.buffer_full_in , 
        \node_1.buffer_full_out , \node_1.receiving_data , 
        \node_1.sending_data , \node_1.data_in , \node_1.data_out , 
        \node_2.clk , \node_2.buffer_full_in , \node_2.buffer_full_out , 
        \node_2.receiving_data , \node_2.sending_data , \node_2.data_in , 
        \node_2.data_out , \node_3.clk , \node_3.buffer_full_in , 
        \node_3.buffer_full_out , \node_3.receiving_data , 
        \node_3.sending_data , \node_3.data_in , \node_3.data_out  );
  input [15:0] \local_node.data_in ;
  output [15:0] \local_node.data_out ;
  input [15:0] \node_0.data_in ;
  output [15:0] \node_0.data_out ;
  input [15:0] \node_1.data_in ;
  output [15:0] \node_1.data_out ;
  input [15:0] \node_2.data_in ;
  output [15:0] \node_2.data_out ;
  input [15:0] \node_3.data_in ;
  output [15:0] \node_3.data_out ;
  input \clk.clk , \reset.reset , \local_node.buffer_full_in ,
         \local_node.receiving_data , \node_0.buffer_full_in ,
         \node_0.receiving_data , \node_1.buffer_full_in ,
         \node_1.receiving_data , \node_2.buffer_full_in ,
         \node_2.receiving_data , \node_3.buffer_full_in ,
         \node_3.receiving_data ;
  output \local_node.buffer_full_out , \local_node.sending_data ,
         \node_0.buffer_full_out , \node_0.sending_data ,
         \node_1.buffer_full_out , \node_1.sending_data ,
         \node_2.buffer_full_out , \node_2.sending_data ,
         \node_3.buffer_full_out , \node_3.sending_data ;
  inout \local_node.clk ,  \node_0.clk ,  \node_1.clk ,  \node_2.clk , 
     \node_3.clk ;
  wire   \buffer_out[4][15] , \buffer_out[4][14] , \buffer_out[4][13] ,
         \buffer_out[4][12] , \buffer_out[4][11] , \buffer_out[4][10] ,
         \buffer_out[4][9] , \buffer_out[4][8] , \buffer_out[4][7] ,
         \buffer_out[4][6] , \buffer_out[4][5] , \buffer_out[4][4] ,
         \buffer_out[4][3] , \buffer_out[4][2] , \buffer_out[4][1] ,
         \buffer_out[4][0] , \buffer_out[3][15] , \buffer_out[3][14] ,
         \buffer_out[3][13] , \buffer_out[3][12] , \buffer_out[3][11] ,
         \buffer_out[3][10] , \buffer_out[3][9] , \buffer_out[3][8] ,
         \buffer_out[3][7] , \buffer_out[3][6] , \buffer_out[3][5] ,
         \buffer_out[3][4] , \buffer_out[3][3] , \buffer_out[3][2] ,
         \buffer_out[3][1] , \buffer_out[3][0] , \buffer_out[2][15] ,
         \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] ,
         \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] ,
         \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] ,
         \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] ,
         \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] ,
         \buffer_out[1][15] , \buffer_out[1][14] , \buffer_out[1][13] ,
         \buffer_out[1][12] , \buffer_out[1][11] , \buffer_out[1][10] ,
         \buffer_out[1][9] , \buffer_out[1][8] , \buffer_out[1][7] ,
         \buffer_out[1][6] , \buffer_out[1][5] , \buffer_out[1][4] ,
         \buffer_out[1][3] , \buffer_out[1][2] , \buffer_out[1][1] ,
         \buffer_out[1][0] , \buffer_out[0][15] , \buffer_out[0][14] ,
         \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] ,
         \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] ,
         \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] ,
         \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] ,
         \buffer_out[0][1] , \buffer_out[0][0] , \next_buffer_out[4][15] ,
         \next_buffer_out[4][14] , \next_buffer_out[4][13] ,
         \next_buffer_out[4][12] , \next_buffer_out[4][11] ,
         \next_buffer_out[4][10] , \next_buffer_out[4][9] ,
         \next_buffer_out[4][8] , \next_buffer_out[4][7] ,
         \next_buffer_out[4][6] , \next_buffer_out[4][5] ,
         \next_buffer_out[4][4] , \next_buffer_out[4][3] ,
         \next_buffer_out[4][2] , \next_buffer_out[4][1] ,
         \next_buffer_out[4][0] , \next_buffer_out[3][15] ,
         \next_buffer_out[3][14] , \next_buffer_out[3][13] ,
         \next_buffer_out[3][12] , \next_buffer_out[3][11] ,
         \next_buffer_out[3][10] , \next_buffer_out[3][9] ,
         \next_buffer_out[3][8] , \next_buffer_out[3][7] ,
         \next_buffer_out[3][6] , \next_buffer_out[3][5] ,
         \next_buffer_out[3][4] , \next_buffer_out[3][3] ,
         \next_buffer_out[3][2] , \next_buffer_out[3][1] ,
         \next_buffer_out[3][0] , \next_buffer_out[2][15] ,
         \next_buffer_out[2][14] , \next_buffer_out[2][13] ,
         \next_buffer_out[2][12] , \next_buffer_out[2][11] ,
         \next_buffer_out[2][10] , \next_buffer_out[2][9] ,
         \next_buffer_out[2][8] , \next_buffer_out[2][7] ,
         \next_buffer_out[2][6] , \next_buffer_out[2][5] ,
         \next_buffer_out[2][4] , \next_buffer_out[2][3] ,
         \next_buffer_out[2][2] , \next_buffer_out[2][1] ,
         \next_buffer_out[2][0] , \next_buffer_out[1][15] ,
         \next_buffer_out[1][14] , \next_buffer_out[1][13] ,
         \next_buffer_out[1][12] , \next_buffer_out[1][11] ,
         \next_buffer_out[1][10] , \next_buffer_out[1][9] ,
         \next_buffer_out[1][8] , \next_buffer_out[1][7] ,
         \next_buffer_out[1][6] , \next_buffer_out[1][5] ,
         \next_buffer_out[1][4] , \next_buffer_out[1][3] ,
         \next_buffer_out[1][2] , \next_buffer_out[1][1] ,
         \next_buffer_out[1][0] , \next_buffer_out[0][15] ,
         \next_buffer_out[0][14] , \next_buffer_out[0][13] ,
         \next_buffer_out[0][12] , \next_buffer_out[0][11] ,
         \next_buffer_out[0][10] , \next_buffer_out[0][9] ,
         \next_buffer_out[0][8] , \next_buffer_out[0][7] ,
         \next_buffer_out[0][6] , \next_buffer_out[0][5] ,
         \next_buffer_out[0][4] , \next_buffer_out[0][3] ,
         \next_buffer_out[0][2] , \next_buffer_out[0][1] ,
         \next_buffer_out[0][0] ;
  wire   [4:0] buffer_full_in;
  wire   [4:0] receiving_data;
  wire   [4:0] pop_v;
  wire   [4:0] data_valid;
  wire   [4:0] next_data_valid;
  wire   [1:0] grant_0;
  wire   [1:0] grant_1;
  wire   [3:0] grant_2;
  wire   [3:0] grant_3;
  wire   [3:0] grant_4;
  tri   \local_node.buffer_full_in ;
  tri   \local_node.buffer_full_out ;
  tri   \local_node.receiving_data ;
  tri   \local_node.sending_data ;
  tri   [15:0] \local_node.data_in ;
  tri   [15:0] \local_node.data_out ;

  converter_in_I_n_node_interface_dut__5 c0 ( .\n.buffer_full_in (
        \node_0.buffer_full_in ), .\n.receiving_data (\node_0.receiving_data ), 
        .\n.data_in (\node_0.data_in ), .\n.buffer_full_out (
        \node_0.buffer_full_out ), .\n.sending_data (\node_0.sending_data ), 
        .\n.data_out (\node_0.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_out_I_n_node_interface_dut_ c1 ( .\n.buffer_full_in (
        \node_1.buffer_full_in ), .\n.receiving_data (\node_1.receiving_data ), 
        .\n.data_in (\node_1.data_in ), .\n.buffer_full_out (
        \node_1.buffer_full_out ), .\n.sending_data (\node_1.sending_data ), 
        .\n.data_out (\node_1.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_in_I_n_node_interface_dut__4 c2 ( .\n.buffer_full_in (
        \node_2.buffer_full_in ), .\n.receiving_data (\node_2.receiving_data ), 
        .\n.data_in (\node_2.data_in ), .\n.buffer_full_out (
        \node_2.buffer_full_out ), .\n.sending_data (\node_2.sending_data ), 
        .\n.data_out (\node_2.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_out_I_n_node_interface_dut_ c3 ( .\n.buffer_full_in (
        \node_3.buffer_full_in ), .\n.receiving_data (\node_3.receiving_data ), 
        .\n.data_in (\node_3.data_in ), .\n.buffer_full_out (
        \node_3.buffer_full_out ), .\n.sending_data (\node_3.sending_data ), 
        .\n.data_out (\node_3.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_out_I_n_node_interface_dut_ c4 ( .\n.buffer_full_in (
        \local_node.buffer_full_in ), .\n.receiving_data (
        \local_node.receiving_data ), .\n.data_in (\local_node.data_in ), 
        .\n.buffer_full_out (\local_node.buffer_full_out ), .\n.sending_data (
        \local_node.sending_data ), .\n.data_out (\local_node.data_out ), 
        .buffer_full_in(1'b0), .receiving_data(1'b0), .data_in({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  fifo_kev_14 \genblk1[0].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[0]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[0]), .data_out({\buffer_out[0][15] , 
        \buffer_out[0][14] , \buffer_out[0][13] , \buffer_out[0][12] , 
        \buffer_out[0][11] , \buffer_out[0][10] , \buffer_out[0][9] , 
        \buffer_out[0][8] , \buffer_out[0][7] , \buffer_out[0][6] , 
        \buffer_out[0][5] , \buffer_out[0][4] , \buffer_out[0][3] , 
        \buffer_out[0][2] , \buffer_out[0][1] , \buffer_out[0][0] }), 
        .next_data_out({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] , 
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .next_data_valid(
        next_data_valid[0]) );
  address_counter_14 \genblk1[0].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] }), 
        .buffer_data_valid(next_data_valid[0]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .buffer_pop(
        pop_v[0]), .receiving_data(1'b0) );
  fifo_kev_13 \genblk1[1].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[1]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[1]), .data_out({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), 
        .next_data_out({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] , 
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .next_data_valid(
        next_data_valid[1]) );
  address_counter_13 \genblk1[1].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] }), 
        .buffer_data_valid(next_data_valid[1]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .buffer_pop(
        pop_v[1]), .receiving_data(1'b0) );
  fifo_kev_12 \genblk1[2].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[2]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[2]), .data_out({\buffer_out[2][15] , 
        \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] , 
        \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] , 
        \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] , 
        \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] , 
        \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] }), 
        .next_data_out({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] , 
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .next_data_valid(
        next_data_valid[2]) );
  address_counter_12 \genblk1[2].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] }), 
        .buffer_data_valid(next_data_valid[2]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .buffer_pop(
        pop_v[2]), .receiving_data(1'b0) );
  fifo_kev_11 \genblk1[3].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[3]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[3]), .data_out({\buffer_out[3][15] , 
        \buffer_out[3][14] , \buffer_out[3][13] , \buffer_out[3][12] , 
        \buffer_out[3][11] , \buffer_out[3][10] , \buffer_out[3][9] , 
        \buffer_out[3][8] , \buffer_out[3][7] , \buffer_out[3][6] , 
        \buffer_out[3][5] , \buffer_out[3][4] , \buffer_out[3][3] , 
        \buffer_out[3][2] , \buffer_out[3][1] , \buffer_out[3][0] }), 
        .next_data_out({\next_buffer_out[3][15] , \next_buffer_out[3][14] , 
        \next_buffer_out[3][13] , \next_buffer_out[3][12] , 
        \next_buffer_out[3][11] , \next_buffer_out[3][10] , 
        \next_buffer_out[3][9] , \next_buffer_out[3][8] , 
        \next_buffer_out[3][7] , \next_buffer_out[3][6] , 
        \next_buffer_out[3][5] , \next_buffer_out[3][4] , 
        \next_buffer_out[3][3] , \next_buffer_out[3][2] , 
        \next_buffer_out[3][1] , \next_buffer_out[3][0] }), .next_data_valid(
        next_data_valid[3]) );
  address_counter_11 \genblk1[3].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[3][15] , \next_buffer_out[3][14] , 
        \next_buffer_out[3][13] , \next_buffer_out[3][12] , 
        \next_buffer_out[3][11] , \next_buffer_out[3][10] , 
        \next_buffer_out[3][9] , \next_buffer_out[3][8] }), 
        .buffer_data_valid(next_data_valid[3]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[3][7] , \next_buffer_out[3][6] , 
        \next_buffer_out[3][5] , \next_buffer_out[3][4] , 
        \next_buffer_out[3][3] , \next_buffer_out[3][2] , 
        \next_buffer_out[3][1] , \next_buffer_out[3][0] }), .buffer_pop(
        pop_v[3]), .receiving_data(1'b0) );
  fifo_kev_10 \genblk1[4].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[4]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[4]), .data_out({\buffer_out[4][15] , 
        \buffer_out[4][14] , \buffer_out[4][13] , \buffer_out[4][12] , 
        \buffer_out[4][11] , \buffer_out[4][10] , \buffer_out[4][9] , 
        \buffer_out[4][8] , \buffer_out[4][7] , \buffer_out[4][6] , 
        \buffer_out[4][5] , \buffer_out[4][4] , \buffer_out[4][3] , 
        \buffer_out[4][2] , \buffer_out[4][1] , \buffer_out[4][0] }), 
        .next_data_out({\next_buffer_out[4][15] , \next_buffer_out[4][14] , 
        \next_buffer_out[4][13] , \next_buffer_out[4][12] , 
        \next_buffer_out[4][11] , \next_buffer_out[4][10] , 
        \next_buffer_out[4][9] , \next_buffer_out[4][8] , 
        \next_buffer_out[4][7] , \next_buffer_out[4][6] , 
        \next_buffer_out[4][5] , \next_buffer_out[4][4] , 
        \next_buffer_out[4][3] , \next_buffer_out[4][2] , 
        \next_buffer_out[4][1] , \next_buffer_out[4][0] }), .next_data_valid(
        next_data_valid[4]) );
  address_counter_10 \genblk1[4].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[4][15] , \next_buffer_out[4][14] , 
        \next_buffer_out[4][13] , \next_buffer_out[4][12] , 
        \next_buffer_out[4][11] , \next_buffer_out[4][10] , 
        \next_buffer_out[4][9] , \next_buffer_out[4][8] }), 
        .buffer_data_valid(next_data_valid[4]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[4][7] , \next_buffer_out[4][6] , 
        \next_buffer_out[4][5] , \next_buffer_out[4][4] , 
        \next_buffer_out[4][3] , \next_buffer_out[4][2] , 
        \next_buffer_out[4][1] , \next_buffer_out[4][0] }), .buffer_pop(
        pop_v[4]), .receiving_data(1'b0) );
  controller5_2 ctrl5 ( .clk(\clk.clk ), .rst(\reset.reset ), .packet_addr({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .local_addr({1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 
        1'b0, 1'b1, 1'b0}), .packet_valid(data_valid), .buffer_full_in({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .grant_0(grant_0), .grant_1(grant_1), 
        .grant_2(grant_2), .grant_3(grant_3), .grant_4(grant_4), .pop_v(pop_v)
         );
  mux2_1_5 mux_n ( .data0({\buffer_out[1][15] , \buffer_out[1][14] , 
        \buffer_out[1][13] , \buffer_out[1][12] , \buffer_out[1][11] , 
        \buffer_out[1][10] , \buffer_out[1][9] , \buffer_out[1][8] , 
        \buffer_out[1][7] , \buffer_out[1][6] , \buffer_out[1][5] , 
        \buffer_out[1][4] , \buffer_out[1][3] , \buffer_out[1][2] , 
        \buffer_out[1][1] , \buffer_out[1][0] }), .data1({\buffer_out[4][15] , 
        \buffer_out[4][14] , \buffer_out[4][13] , \buffer_out[4][12] , 
        \buffer_out[4][11] , \buffer_out[4][10] , \buffer_out[4][9] , 
        \buffer_out[4][8] , \buffer_out[4][7] , \buffer_out[4][6] , 
        \buffer_out[4][5] , \buffer_out[4][4] , \buffer_out[4][3] , 
        \buffer_out[4][2] , \buffer_out[4][1] , \buffer_out[4][0] }), 
        .select0(grant_0[0]), .select1(grant_0[1]) );
  mux2_1_4 mux_s ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[4][15] , 
        \buffer_out[4][14] , \buffer_out[4][13] , \buffer_out[4][12] , 
        \buffer_out[4][11] , \buffer_out[4][10] , \buffer_out[4][9] , 
        \buffer_out[4][8] , \buffer_out[4][7] , \buffer_out[4][6] , 
        \buffer_out[4][5] , \buffer_out[4][4] , \buffer_out[4][3] , 
        \buffer_out[4][2] , \buffer_out[4][1] , \buffer_out[4][0] }), 
        .select0(grant_1[0]), .select1(grant_1[1]) );
  mux4_1_8 mux_e ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[3][15] , \buffer_out[3][14] , \buffer_out[3][13] , 
        \buffer_out[3][12] , \buffer_out[3][11] , \buffer_out[3][10] , 
        \buffer_out[3][9] , \buffer_out[3][8] , \buffer_out[3][7] , 
        \buffer_out[3][6] , \buffer_out[3][5] , \buffer_out[3][4] , 
        \buffer_out[3][3] , \buffer_out[3][2] , \buffer_out[3][1] , 
        \buffer_out[3][0] }), .data3({\buffer_out[4][15] , \buffer_out[4][14] , 
        \buffer_out[4][13] , \buffer_out[4][12] , \buffer_out[4][11] , 
        \buffer_out[4][10] , \buffer_out[4][9] , \buffer_out[4][8] , 
        \buffer_out[4][7] , \buffer_out[4][6] , \buffer_out[4][5] , 
        \buffer_out[4][4] , \buffer_out[4][3] , \buffer_out[4][2] , 
        \buffer_out[4][1] , \buffer_out[4][0] }), .select0(grant_2[0]), 
        .select1(grant_2[1]), .select2(grant_2[2]), .select3(grant_2[3]) );
  mux4_1_7 mux_w ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[2][15] , \buffer_out[2][14] , \buffer_out[2][13] , 
        \buffer_out[2][12] , \buffer_out[2][11] , \buffer_out[2][10] , 
        \buffer_out[2][9] , \buffer_out[2][8] , \buffer_out[2][7] , 
        \buffer_out[2][6] , \buffer_out[2][5] , \buffer_out[2][4] , 
        \buffer_out[2][3] , \buffer_out[2][2] , \buffer_out[2][1] , 
        \buffer_out[2][0] }), .data3({\buffer_out[4][15] , \buffer_out[4][14] , 
        \buffer_out[4][13] , \buffer_out[4][12] , \buffer_out[4][11] , 
        \buffer_out[4][10] , \buffer_out[4][9] , \buffer_out[4][8] , 
        \buffer_out[4][7] , \buffer_out[4][6] , \buffer_out[4][5] , 
        \buffer_out[4][4] , \buffer_out[4][3] , \buffer_out[4][2] , 
        \buffer_out[4][1] , \buffer_out[4][0] }), .select0(grant_3[0]), 
        .select1(grant_3[1]), .select2(grant_3[2]), .select3(grant_3[3]) );
  mux4_1_6 mux_l ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[2][15] , \buffer_out[2][14] , \buffer_out[2][13] , 
        \buffer_out[2][12] , \buffer_out[2][11] , \buffer_out[2][10] , 
        \buffer_out[2][9] , \buffer_out[2][8] , \buffer_out[2][7] , 
        \buffer_out[2][6] , \buffer_out[2][5] , \buffer_out[2][4] , 
        \buffer_out[2][3] , \buffer_out[2][2] , \buffer_out[2][1] , 
        \buffer_out[2][0] }), .data3({\buffer_out[3][15] , \buffer_out[3][14] , 
        \buffer_out[3][13] , \buffer_out[3][12] , \buffer_out[3][11] , 
        \buffer_out[3][10] , \buffer_out[3][9] , \buffer_out[3][8] , 
        \buffer_out[3][7] , \buffer_out[3][6] , \buffer_out[3][5] , 
        \buffer_out[3][4] , \buffer_out[3][3] , \buffer_out[3][2] , 
        \buffer_out[3][1] , \buffer_out[3][0] }), .select0(grant_4[0]), 
        .select1(grant_4[1]), .select2(grant_4[2]), .select3(grant_4[3]) );
endmodule


module converter_in_I_n_node_interface_dut__3 ( \n.buffer_full_in , 
        \n.receiving_data , \n.data_in , \n.buffer_full_out , \n.sending_data , 
        \n.data_out , buffer_full_out, sending_data, data_out, buffer_full_in, 
        receiving_data, data_in );
  input [15:0] \n.data_in ;
  output [15:0] \n.data_out ;
  output [15:0] data_out;
  input [15:0] data_in;
  input \n.buffer_full_in , \n.receiving_data , buffer_full_in, receiving_data;
  output \n.buffer_full_out , \n.sending_data , buffer_full_out, sending_data;
  wire   \n.buffer_full_in , \n.receiving_data , buffer_full_in,
         receiving_data;
  assign buffer_full_out = \n.buffer_full_in ;
  assign sending_data = \n.receiving_data ;
  assign data_out[15] = \n.data_in  [15];
  assign data_out[14] = \n.data_in  [14];
  assign data_out[13] = \n.data_in  [13];
  assign data_out[12] = \n.data_in  [12];
  assign data_out[11] = \n.data_in  [11];
  assign data_out[10] = \n.data_in  [10];
  assign data_out[9] = \n.data_in  [9];
  assign data_out[8] = \n.data_in  [8];
  assign data_out[7] = \n.data_in  [7];
  assign data_out[6] = \n.data_in  [6];
  assign data_out[5] = \n.data_in  [5];
  assign data_out[4] = \n.data_in  [4];
  assign data_out[3] = \n.data_in  [3];
  assign data_out[2] = \n.data_in  [2];
  assign data_out[1] = \n.data_in  [1];
  assign data_out[0] = \n.data_in  [0];
  assign \n.buffer_full_out  = buffer_full_in;
  assign \n.sending_data  = receiving_data;
  assign \n.data_out  [15] = data_in[15];
  assign \n.data_out  [14] = data_in[14];
  assign \n.data_out  [13] = data_in[13];
  assign \n.data_out  [12] = data_in[12];
  assign \n.data_out  [11] = data_in[11];
  assign \n.data_out  [10] = data_in[10];
  assign \n.data_out  [9] = data_in[9];
  assign \n.data_out  [8] = data_in[8];
  assign \n.data_out  [7] = data_in[7];
  assign \n.data_out  [6] = data_in[6];
  assign \n.data_out  [5] = data_in[5];
  assign \n.data_out  [4] = data_in[4];
  assign \n.data_out  [3] = data_in[3];
  assign \n.data_out  [2] = data_in[2];
  assign \n.data_out  [1] = data_in[1];
  assign \n.data_out  [0] = data_in[0];

endmodule


module converter_in_I_n_node_interface_dut__2 ( \n.buffer_full_in , 
        \n.receiving_data , \n.data_in , \n.buffer_full_out , \n.sending_data , 
        \n.data_out , buffer_full_out, sending_data, data_out, buffer_full_in, 
        receiving_data, data_in );
  input [15:0] \n.data_in ;
  output [15:0] \n.data_out ;
  output [15:0] data_out;
  input [15:0] data_in;
  input \n.buffer_full_in , \n.receiving_data , buffer_full_in, receiving_data;
  output \n.buffer_full_out , \n.sending_data , buffer_full_out, sending_data;
  wire   \n.buffer_full_in , \n.receiving_data , buffer_full_in,
         receiving_data;
  assign buffer_full_out = \n.buffer_full_in ;
  assign sending_data = \n.receiving_data ;
  assign data_out[15] = \n.data_in  [15];
  assign data_out[14] = \n.data_in  [14];
  assign data_out[13] = \n.data_in  [13];
  assign data_out[12] = \n.data_in  [12];
  assign data_out[11] = \n.data_in  [11];
  assign data_out[10] = \n.data_in  [10];
  assign data_out[9] = \n.data_in  [9];
  assign data_out[8] = \n.data_in  [8];
  assign data_out[7] = \n.data_in  [7];
  assign data_out[6] = \n.data_in  [6];
  assign data_out[5] = \n.data_in  [5];
  assign data_out[4] = \n.data_in  [4];
  assign data_out[3] = \n.data_in  [3];
  assign data_out[2] = \n.data_in  [2];
  assign data_out[1] = \n.data_in  [1];
  assign data_out[0] = \n.data_in  [0];
  assign \n.buffer_full_out  = buffer_full_in;
  assign \n.sending_data  = receiving_data;
  assign \n.data_out  [15] = data_in[15];
  assign \n.data_out  [14] = data_in[14];
  assign \n.data_out  [13] = data_in[13];
  assign \n.data_out  [12] = data_in[12];
  assign \n.data_out  [11] = data_in[11];
  assign \n.data_out  [10] = data_in[10];
  assign \n.data_out  [9] = data_in[9];
  assign \n.data_out  [8] = data_in[8];
  assign \n.data_out  [7] = data_in[7];
  assign \n.data_out  [6] = data_in[6];
  assign \n.data_out  [5] = data_in[5];
  assign \n.data_out  [4] = data_in[4];
  assign \n.data_out  [3] = data_in[3];
  assign \n.data_out  [2] = data_in[2];
  assign \n.data_out  [1] = data_in[1];
  assign \n.data_out  [0] = data_in[0];

endmodule


module fifo_kev_9 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_19 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_9 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_19 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_18 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_9 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_18 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_9_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_9 ( clk, rst, interface_flit_length, buffer_flit_length, 
        buffer_data_valid, interface_flit_address, buffer_flit_address, 
        buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_9 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_9 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_9_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), .SUM(
        {SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_8 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_17 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_8 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_17 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_16 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_8 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_16 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_8_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_8 ( clk, rst, interface_flit_length, buffer_flit_length, 
        buffer_data_valid, interface_flit_address, buffer_flit_address, 
        buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_8 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_8 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_8_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), .SUM(
        {SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_7 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_15 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_7 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_15 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_14 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_7 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_14 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_7_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_7 ( clk, rst, interface_flit_length, buffer_flit_length, 
        buffer_data_valid, interface_flit_address, buffer_flit_address, 
        buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_7 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_7 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_7_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), .SUM(
        {SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_6 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_13 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_6 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_13 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_12 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_6 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_12 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_6_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_6 ( clk, rst, interface_flit_length, buffer_flit_length, 
        buffer_data_valid, interface_flit_address, buffer_flit_address, 
        buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_6 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_6 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_6_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), .SUM(
        {SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_5 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_11 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_5 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_11 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_10 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_5 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_10 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, 
        n15, n13, n11, n9, n7, n5}) );
endmodule


module address_counter_5_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_5 ( clk, rst, interface_flit_length, buffer_flit_length, 
        buffer_data_valid, interface_flit_address, buffer_flit_address, 
        buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_5 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_5 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_5_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), .SUM(
        {SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module flipflop_BITS2_3 ( clk, data_i, data_o );
  input [1:0] data_i;
  output [1:0] data_o;
  input clk;


  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS2_3 ( clk, enable_i, reset, data_i, data_o );
  input [1:0] data_i;
  input [1:0] data_o;
  input clk, enable_i, reset;
  wire   n10, n11, n1, n5, n7, n8, n9;
  wire   [1:0] write_data;

  AOI22X1 U5 ( .IN1(enable_i), .IN2(data_i[1]), .IN3(n10), .IN4(n1), .QN(n9)
         );
  AOI22X1 U6 ( .IN1(data_i[0]), .IN2(enable_i), .IN3(n11), .IN4(n1), .QN(n8)
         );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n9), .QN(write_data[1]) );
  NOR2X0 U4 ( .IN1(reset), .IN2(n8), .QN(write_data[0]) );
  AND2X1 U7 ( .IN1(data_o[1]), .IN2(n7), .Q(n10) );
  AND2X1 U8 ( .IN1(data_o[0]), .IN2(n5), .Q(n11) );
  flipflop_BITS2_3 FF ( .clk(clk), .data_i(write_data), .data_o({n7, n5}) );
endmodule


module flipflop_BITS1_15 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_15 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_15 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter2_3 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [1:0] request;
  output [1:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   tail_en, n1, n2;
  wire   [1:0] req_i;
  wire   [1:0] req_o;

  AND3X1 U10 ( .IN1(request[1]), .IN2(n1), .IN3(n2), .Q(grant[1]) );
  AND3X1 U11 ( .IN1(request[0]), .IN2(n2), .IN3(request[1]), .Q(tail_en) );
  INVX0 U6 ( .INP(request[0]), .ZN(n1) );
  NOR2X0 U7 ( .IN1(buffer_full_i), .IN2(n1), .QN(grant[0]) );
  INVX0 U8 ( .INP(buffer_full_i), .ZN(n2) );
  OA21X1 U9 ( .IN1(request[1]), .IN2(request[0]), .IN3(n2), .Q(grant_v_o) );
  register_BITS2_3 req_record ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i({1'b1, 1'b0}), .data_o({1'b0, 1'b0}) );
  register_BITS1_15 tail ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i(1'b1), .data_o(1'b0) );
endmodule


module flipflop_BITS2_2 ( clk, data_i, data_o );
  input [1:0] data_i;
  output [1:0] data_o;
  input clk;


  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS2_2 ( clk, enable_i, reset, data_i, data_o );
  input [1:0] data_i;
  input [1:0] data_o;
  input clk, enable_i, reset;
  wire   n10, n11, n1, n5, n7, n8, n9;
  wire   [1:0] write_data;

  AOI22X1 U5 ( .IN1(enable_i), .IN2(data_i[1]), .IN3(n10), .IN4(n1), .QN(n9)
         );
  AOI22X1 U6 ( .IN1(data_i[0]), .IN2(enable_i), .IN3(n11), .IN4(n1), .QN(n8)
         );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n9), .QN(write_data[1]) );
  NOR2X0 U4 ( .IN1(reset), .IN2(n8), .QN(write_data[0]) );
  AND2X1 U7 ( .IN1(data_o[1]), .IN2(n7), .Q(n10) );
  AND2X1 U8 ( .IN1(data_o[0]), .IN2(n5), .Q(n11) );
  flipflop_BITS2_2 FF ( .clk(clk), .data_i(write_data), .data_o({n7, n5}) );
endmodule


module flipflop_BITS1_14 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_14 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_14 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter2_2 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [1:0] request;
  output [1:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   tail_en, n1, n2;
  wire   [1:0] req_i;
  wire   [1:0] req_o;

  AND3X1 U10 ( .IN1(request[1]), .IN2(n1), .IN3(n2), .Q(grant[1]) );
  AND3X1 U11 ( .IN1(request[0]), .IN2(n2), .IN3(request[1]), .Q(tail_en) );
  INVX0 U6 ( .INP(request[0]), .ZN(n1) );
  NOR2X0 U7 ( .IN1(buffer_full_i), .IN2(n1), .QN(grant[0]) );
  INVX0 U8 ( .INP(buffer_full_i), .ZN(n2) );
  OA21X1 U9 ( .IN1(request[1]), .IN2(request[0]), .IN3(n2), .Q(grant_v_o) );
  register_BITS2_2 req_record ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i({1'b1, 1'b0}), .data_o({1'b0, 1'b0}) );
  register_BITS1_14 tail ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i(1'b1), .data_o(1'b0) );
endmodule


module flipflop_BITS4_17 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_17 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_17 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS4_16 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_16 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_16 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS4_15 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_15 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_15 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS1_13 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_13 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_13 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_12 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_12 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_12 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter4_5 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [3:0] request;
  output [3:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[2][3] , \req_i[2][2] , \req_i[2][1] , \req_i[2][0] ,
         \req_i[1][3] , \req_i[1][2] , \req_i[1][1] , \req_i[1][0] ,
         \req_i[0][3] , \req_i[0][2] , \req_i[0][1] , tail_en, N71, N265, N266,
         N267, N268, N276, N282, N291, N300, N301, N302, N303, n1, n2, n3, n4,
         n6, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21;
  wire   [2:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N265 = request[0];
  assign N266 = request[1];
  assign N267 = request[2];
  assign N268 = request[3];

  LATCHX1 shift_reg ( .CLK(1'b0), .D(1'b0), .Q(N71) );
  LATCHX1 \grant_reg[3]  ( .CLK(1'b1), .D(N303), .Q(grant[3]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N302), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N301), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N300), .Q(grant[0]) );
  LNANDX1 \req_i_reg[2][3]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][3] ) );
  LNANDX1 \req_i_reg[2][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][2] ) );
  LNANDX1 \req_i_reg[2][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][1] ) );
  LNANDX1 \req_i_reg[2][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][0] ) );
  LNANDX1 \req_i_reg[1][3]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][3] ) );
  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][3]  ( .CLK(tail_en), .D(N282), .Q(\req_i[0][3] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(n1), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(n4), .Q(\req_i[0][1] ) );
  LATCHX1 \tail_i_reg[0]  ( .CLK(tail_en), .D(N276), .Q(tail_i[0]) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N291), .D(tail_en), .Q(req_en[0]) );
  AND3X1 U35 ( .IN1(grant_v_o), .IN2(n19), .IN3(N267), .Q(N302) );
  NAND4X0 U37 ( .IN1(n17), .IN2(grant_v_o), .IN3(n16), .IN4(n20), .QN(N291) );
  AO21X1 U38 ( .IN1(n14), .IN2(n19), .IN3(buffer_full_i), .Q(n21) );
  NOR3X0 U39 ( .IN1(n4), .IN2(N282), .IN3(n1), .QN(n17) );
  NAND4X0 U41 ( .IN1(n11), .IN2(n13), .IN3(n9), .IN4(n10), .QN(N276) );
  AOI22X1 U42 ( .IN1(n2), .IN2(n15), .IN3(n15), .IN4(N265), .QN(n13) );
  AND2X1 U43 ( .IN1(N268), .IN2(n6), .Q(n15) );
  OA22X1 U44 ( .IN1(n6), .IN2(n18), .IN3(n6), .IN4(n3), .Q(n11) );
  INVX0 U15 ( .INP(N267), .ZN(n6) );
  INVX0 U16 ( .INP(n18), .ZN(n2) );
  NAND2X1 U17 ( .IN1(N266), .IN2(N265), .QN(n10) );
  NAND2X1 U18 ( .IN1(N267), .IN2(N268), .QN(n12) );
  INVX0 U19 ( .INP(N265), .ZN(n3) );
  NAND2X1 U20 ( .IN1(N266), .IN2(n3), .QN(n18) );
  NOR2X0 U21 ( .IN1(N266), .IN2(N265), .QN(n19) );
  INVX0 U22 ( .INP(n21), .ZN(grant_v_o) );
  NOR2X0 U23 ( .IN1(N268), .IN2(N267), .QN(n14) );
  NAND2X1 U24 ( .IN1(n15), .IN2(n19), .QN(n20) );
  NOR2X0 U25 ( .IN1(N265), .IN2(n2), .QN(n16) );
  NAND2X1 U26 ( .IN1(N71), .IN2(n7), .QN(n9) );
  INVX0 U27 ( .INP(n12), .ZN(n7) );
  INVX0 U28 ( .INP(n10), .ZN(n4) );
  INVX0 U29 ( .INP(n11), .ZN(n1) );
  NAND2X1 U30 ( .IN1(n13), .IN2(n12), .QN(N282) );
  NOR2X0 U31 ( .IN1(n21), .IN2(n17), .QN(tail_en) );
  NOR2X0 U32 ( .IN1(n3), .IN2(n21), .QN(N300) );
  NOR2X0 U33 ( .IN1(n18), .IN2(n21), .QN(N301) );
  NOR2X0 U34 ( .IN1(n21), .IN2(n20), .QN(N303) );
  register_BITS4_17 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][3] , \req_i[0][2] , \req_i[0][1] , 
        1'b0}), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS4_16 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][3] , \req_i[1][2] , \req_i[1][1] , 
        \req_i[1][0] }), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS4_15 \genblk1[2].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[2][3] , \req_i[2][2] , \req_i[2][1] , 
        \req_i[2][0] }), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS1_13 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(tail_i[0]), .data_o(1'b0) );
  register_BITS1_12 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module flipflop_BITS4_14 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_14 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_14 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS4_13 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_13 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_13 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS4_12 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_12 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_12 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS1_11 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_11 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_11 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_10 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_10 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_10 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter4_4 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [3:0] request;
  output [3:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[2][3] , \req_i[2][2] , \req_i[2][1] , \req_i[2][0] ,
         \req_i[1][3] , \req_i[1][2] , \req_i[1][1] , \req_i[1][0] ,
         \req_i[0][3] , \req_i[0][2] , \req_i[0][1] , tail_en, N71, N265, N266,
         N267, N268, N276, N282, N291, N300, N301, N302, N303, n1, n2, n3, n4,
         n6, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21;
  wire   [2:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N265 = request[0];
  assign N266 = request[1];
  assign N267 = request[2];
  assign N268 = request[3];

  LATCHX1 shift_reg ( .CLK(1'b0), .D(1'b0), .Q(N71) );
  LATCHX1 \grant_reg[3]  ( .CLK(1'b1), .D(N303), .Q(grant[3]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N302), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N301), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N300), .Q(grant[0]) );
  LNANDX1 \req_i_reg[2][3]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][3] ) );
  LNANDX1 \req_i_reg[2][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][2] ) );
  LNANDX1 \req_i_reg[2][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][1] ) );
  LNANDX1 \req_i_reg[2][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][0] ) );
  LNANDX1 \req_i_reg[1][3]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][3] ) );
  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][3]  ( .CLK(tail_en), .D(N282), .Q(\req_i[0][3] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(n1), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(n4), .Q(\req_i[0][1] ) );
  LATCHX1 \tail_i_reg[0]  ( .CLK(tail_en), .D(N276), .Q(tail_i[0]) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N291), .D(tail_en), .Q(req_en[0]) );
  AND3X1 U35 ( .IN1(grant_v_o), .IN2(n19), .IN3(N267), .Q(N302) );
  NAND4X0 U37 ( .IN1(n17), .IN2(grant_v_o), .IN3(n16), .IN4(n20), .QN(N291) );
  AO21X1 U38 ( .IN1(n14), .IN2(n19), .IN3(buffer_full_i), .Q(n21) );
  NOR3X0 U39 ( .IN1(n4), .IN2(N282), .IN3(n1), .QN(n17) );
  NAND4X0 U41 ( .IN1(n11), .IN2(n13), .IN3(n9), .IN4(n10), .QN(N276) );
  AOI22X1 U42 ( .IN1(n2), .IN2(n15), .IN3(n15), .IN4(N265), .QN(n13) );
  AND2X1 U43 ( .IN1(N268), .IN2(n6), .Q(n15) );
  OA22X1 U44 ( .IN1(n6), .IN2(n18), .IN3(n6), .IN4(n3), .Q(n11) );
  INVX0 U15 ( .INP(N267), .ZN(n6) );
  INVX0 U16 ( .INP(n18), .ZN(n2) );
  NAND2X1 U17 ( .IN1(N266), .IN2(N265), .QN(n10) );
  NAND2X1 U18 ( .IN1(N267), .IN2(N268), .QN(n12) );
  INVX0 U19 ( .INP(N265), .ZN(n3) );
  NAND2X1 U20 ( .IN1(N266), .IN2(n3), .QN(n18) );
  NOR2X0 U21 ( .IN1(N266), .IN2(N265), .QN(n19) );
  INVX0 U22 ( .INP(n21), .ZN(grant_v_o) );
  NOR2X0 U23 ( .IN1(N268), .IN2(N267), .QN(n14) );
  NAND2X1 U24 ( .IN1(n15), .IN2(n19), .QN(n20) );
  NOR2X0 U25 ( .IN1(N265), .IN2(n2), .QN(n16) );
  NAND2X1 U26 ( .IN1(N71), .IN2(n7), .QN(n9) );
  INVX0 U27 ( .INP(n12), .ZN(n7) );
  INVX0 U28 ( .INP(n10), .ZN(n4) );
  INVX0 U29 ( .INP(n11), .ZN(n1) );
  NAND2X1 U30 ( .IN1(n13), .IN2(n12), .QN(N282) );
  NOR2X0 U31 ( .IN1(n21), .IN2(n17), .QN(tail_en) );
  NOR2X0 U32 ( .IN1(n3), .IN2(n21), .QN(N300) );
  NOR2X0 U33 ( .IN1(n18), .IN2(n21), .QN(N301) );
  NOR2X0 U34 ( .IN1(n21), .IN2(n20), .QN(N303) );
  register_BITS4_14 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][3] , \req_i[0][2] , \req_i[0][1] , 
        1'b0}), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS4_13 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][3] , \req_i[1][2] , \req_i[1][1] , 
        \req_i[1][0] }), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS4_12 \genblk1[2].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[2][3] , \req_i[2][2] , \req_i[2][1] , 
        \req_i[2][0] }), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS1_11 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(tail_i[0]), .data_o(1'b0) );
  register_BITS1_10 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module flipflop_BITS4_11 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_11 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_11 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS4_10 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_10 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_10 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS4_9 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_9 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_9 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS1_9 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_9 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_9 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_8 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_8 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_8 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter4_3 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [3:0] request;
  output [3:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[2][3] , \req_i[2][2] , \req_i[2][1] , \req_i[2][0] ,
         \req_i[1][3] , \req_i[1][2] , \req_i[1][1] , \req_i[1][0] ,
         \req_i[0][3] , \req_i[0][2] , \req_i[0][1] , tail_en, N71, N265, N266,
         N267, N268, N276, N282, N291, N300, N301, N302, N303, n1, n2, n3, n4,
         n6, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21;
  wire   [2:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N265 = request[0];
  assign N266 = request[1];
  assign N267 = request[2];
  assign N268 = request[3];

  LATCHX1 shift_reg ( .CLK(1'b0), .D(1'b0), .Q(N71) );
  LATCHX1 \grant_reg[3]  ( .CLK(1'b1), .D(N303), .Q(grant[3]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N302), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N301), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N300), .Q(grant[0]) );
  LNANDX1 \req_i_reg[2][3]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][3] ) );
  LNANDX1 \req_i_reg[2][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][2] ) );
  LNANDX1 \req_i_reg[2][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][1] ) );
  LNANDX1 \req_i_reg[2][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][0] ) );
  LNANDX1 \req_i_reg[1][3]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][3] ) );
  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][3]  ( .CLK(tail_en), .D(N282), .Q(\req_i[0][3] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(n1), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(n4), .Q(\req_i[0][1] ) );
  LATCHX1 \tail_i_reg[0]  ( .CLK(tail_en), .D(N276), .Q(tail_i[0]) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N291), .D(tail_en), .Q(req_en[0]) );
  AND3X1 U35 ( .IN1(grant_v_o), .IN2(n19), .IN3(N267), .Q(N302) );
  NAND4X0 U37 ( .IN1(n17), .IN2(grant_v_o), .IN3(n16), .IN4(n20), .QN(N291) );
  AO21X1 U38 ( .IN1(n14), .IN2(n19), .IN3(buffer_full_i), .Q(n21) );
  NOR3X0 U39 ( .IN1(n4), .IN2(N282), .IN3(n1), .QN(n17) );
  NAND4X0 U41 ( .IN1(n11), .IN2(n13), .IN3(n9), .IN4(n10), .QN(N276) );
  AOI22X1 U42 ( .IN1(n2), .IN2(n15), .IN3(n15), .IN4(N265), .QN(n13) );
  AND2X1 U43 ( .IN1(N268), .IN2(n6), .Q(n15) );
  OA22X1 U44 ( .IN1(n6), .IN2(n18), .IN3(n6), .IN4(n3), .Q(n11) );
  INVX0 U15 ( .INP(N267), .ZN(n6) );
  INVX0 U16 ( .INP(n18), .ZN(n2) );
  NAND2X1 U17 ( .IN1(N266), .IN2(N265), .QN(n10) );
  NAND2X1 U18 ( .IN1(N267), .IN2(N268), .QN(n12) );
  INVX0 U19 ( .INP(N265), .ZN(n3) );
  NAND2X1 U20 ( .IN1(N266), .IN2(n3), .QN(n18) );
  NOR2X0 U21 ( .IN1(N266), .IN2(N265), .QN(n19) );
  INVX0 U22 ( .INP(n21), .ZN(grant_v_o) );
  NOR2X0 U23 ( .IN1(N268), .IN2(N267), .QN(n14) );
  NAND2X1 U24 ( .IN1(n15), .IN2(n19), .QN(n20) );
  NOR2X0 U25 ( .IN1(N265), .IN2(n2), .QN(n16) );
  NAND2X1 U26 ( .IN1(N71), .IN2(n7), .QN(n9) );
  INVX0 U27 ( .INP(n12), .ZN(n7) );
  INVX0 U28 ( .INP(n10), .ZN(n4) );
  INVX0 U29 ( .INP(n11), .ZN(n1) );
  NAND2X1 U30 ( .IN1(n13), .IN2(n12), .QN(N282) );
  NOR2X0 U31 ( .IN1(n21), .IN2(n17), .QN(tail_en) );
  NOR2X0 U32 ( .IN1(n3), .IN2(n21), .QN(N300) );
  NOR2X0 U33 ( .IN1(n18), .IN2(n21), .QN(N301) );
  NOR2X0 U34 ( .IN1(n21), .IN2(n20), .QN(N303) );
  register_BITS4_11 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][3] , \req_i[0][2] , \req_i[0][1] , 
        1'b0}), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS4_10 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][3] , \req_i[1][2] , \req_i[1][1] , 
        \req_i[1][0] }), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS4_9 \genblk1[2].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[2][3] , \req_i[2][2] , \req_i[2][1] , 
        \req_i[2][0] }), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS1_9 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(tail_i[0]), .data_o(1'b0) );
  register_BITS1_8 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module dccl_9 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_8 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_7 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_6 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_5 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module controller5_1 ( clk, rst, .packet_addr({\packet_addr[4][7] , 
        \packet_addr[4][6] , \packet_addr[4][5] , \packet_addr[4][4] , 
        \packet_addr[4][3] , \packet_addr[4][2] , \packet_addr[4][1] , 
        \packet_addr[4][0] , \packet_addr[3][7] , \packet_addr[3][6] , 
        \packet_addr[3][5] , \packet_addr[3][4] , \packet_addr[3][3] , 
        \packet_addr[3][2] , \packet_addr[3][1] , \packet_addr[3][0] , 
        \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] , 
        \packet_addr[2][4] , \packet_addr[2][3] , \packet_addr[2][2] , 
        \packet_addr[2][1] , \packet_addr[2][0] , \packet_addr[1][7] , 
        \packet_addr[1][6] , \packet_addr[1][5] , \packet_addr[1][4] , 
        \packet_addr[1][3] , \packet_addr[1][2] , \packet_addr[1][1] , 
        \packet_addr[1][0] , \packet_addr[0][7] , \packet_addr[0][6] , 
        \packet_addr[0][5] , \packet_addr[0][4] , \packet_addr[0][3] , 
        \packet_addr[0][2] , \packet_addr[0][1] , \packet_addr[0][0] }), 
        local_addr, packet_valid, buffer_full_in, grant_0, grant_1, grant_2, 
        grant_3, grant_4, grant_v, pop_v );
  input [7:0] local_addr;
  input [4:0] packet_valid;
  input [4:0] buffer_full_in;
  output [1:0] grant_0;
  output [1:0] grant_1;
  output [3:0] grant_2;
  output [3:0] grant_3;
  output [3:0] grant_4;
  output [4:0] grant_v;
  output [4:0] pop_v;
  input clk, rst, \packet_addr[4][7] , \packet_addr[4][6] ,
         \packet_addr[4][5] , \packet_addr[4][4] , \packet_addr[4][3] ,
         \packet_addr[4][2] , \packet_addr[4][1] , \packet_addr[4][0] ,
         \packet_addr[3][7] , \packet_addr[3][6] , \packet_addr[3][5] ,
         \packet_addr[3][4] , \packet_addr[3][3] , \packet_addr[3][2] ,
         \packet_addr[3][1] , \packet_addr[3][0] , \packet_addr[2][7] ,
         \packet_addr[2][6] , \packet_addr[2][5] , \packet_addr[2][4] ,
         \packet_addr[2][3] , \packet_addr[2][2] , \packet_addr[2][1] ,
         \packet_addr[2][0] , \packet_addr[1][7] , \packet_addr[1][6] ,
         \packet_addr[1][5] , \packet_addr[1][4] , \packet_addr[1][3] ,
         \packet_addr[1][2] , \packet_addr[1][1] , \packet_addr[1][0] ,
         \packet_addr[0][7] , \packet_addr[0][6] , \packet_addr[0][5] ,
         \packet_addr[0][4] , \packet_addr[0][3] , \packet_addr[0][2] ,
         \packet_addr[0][1] , \packet_addr[0][0] ;
  wire   \request[4][3] , \request[4][2] , \request[4][1] , \request[4][0] ,
         \request[3][3] , \request[3][2] , \request[3][1] , \request[3][0] ,
         \request[2][3] , \request[2][2] , \request[2][1] , \request[2][0] ,
         \request[1][1] , \request[1][0] , \request[0][1] , \request[0][0] ;

  OR4X1 U1 ( .IN1(grant_1[1]), .IN2(grant_0[1]), .IN3(grant_3[3]), .IN4(
        grant_2[3]), .Q(pop_v[4]) );
  OR2X1 U2 ( .IN1(grant_2[2]), .IN2(grant_4[3]), .Q(pop_v[3]) );
  OR2X1 U3 ( .IN1(grant_3[2]), .IN2(grant_4[2]), .Q(pop_v[2]) );
  OR4X1 U4 ( .IN1(grant_2[1]), .IN2(grant_0[0]), .IN3(grant_4[1]), .IN4(
        grant_3[1]), .Q(pop_v[1]) );
  OR4X1 U5 ( .IN1(grant_2[0]), .IN2(grant_1[0]), .IN3(grant_4[0]), .IN4(
        grant_3[0]), .Q(pop_v[0]) );
  arbiter2_3 arbiter_n ( .clk(clk), .rst(rst), .request({\request[0][1] , 
        \request[0][0] }), .buffer_full_i(buffer_full_in[0]), .grant(grant_0), 
        .grant_v_o(grant_v[0]) );
  arbiter2_2 arbiter_s ( .clk(clk), .rst(rst), .request({\request[1][1] , 
        \request[1][0] }), .buffer_full_i(buffer_full_in[1]), .grant(grant_1), 
        .grant_v_o(grant_v[1]) );
  arbiter4_5 arbiter_e ( .clk(clk), .rst(rst), .request({\request[2][3] , 
        \request[2][2] , \request[2][1] , \request[2][0] }), .buffer_full_i(
        buffer_full_in[2]), .grant(grant_2), .grant_v_o(grant_v[2]) );
  arbiter4_4 arbiter_w ( .clk(clk), .rst(rst), .request({\request[3][3] , 
        \request[3][2] , \request[3][1] , \request[3][0] }), .buffer_full_i(
        buffer_full_in[3]), .grant(grant_3), .grant_v_o(grant_v[3]) );
  arbiter4_3 arbiter_l ( .clk(clk), .rst(rst), .request({\request[4][3] , 
        \request[4][2] , \request[4][1] , \request[4][0] }), .buffer_full_i(
        buffer_full_in[4]), .grant(grant_4), .grant_v_o(grant_v[4]) );
  dccl_9 dccl_n ( .packet_addr_y_i({\packet_addr[0][3] , \packet_addr[0][2] , 
        \packet_addr[0][1] , \packet_addr[0][0] }), .packet_addr_x_i({
        \packet_addr[0][7] , \packet_addr[0][6] , \packet_addr[0][5] , 
        \packet_addr[0][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[0]), 
        .east_req(\request[2][0] ), .south_req(\request[1][0] ), .west_req(
        \request[3][0] ), .local_req(\request[4][0] ) );
  dccl_8 dccl_s ( .packet_addr_y_i({\packet_addr[1][3] , \packet_addr[1][2] , 
        \packet_addr[1][1] , \packet_addr[1][0] }), .packet_addr_x_i({
        \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] , 
        \packet_addr[1][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[1]), 
        .north_req(\request[0][0] ), .east_req(\request[2][1] ), .west_req(
        \request[3][1] ), .local_req(\request[4][1] ) );
  dccl_7 dccl_e ( .packet_addr_y_i({\packet_addr[2][3] , \packet_addr[2][2] , 
        \packet_addr[2][1] , \packet_addr[2][0] }), .packet_addr_x_i({
        \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] , 
        \packet_addr[2][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[2]), 
        .west_req(\request[3][2] ), .local_req(\request[4][2] ) );
  dccl_6 dccl_w ( .packet_addr_y_i({\packet_addr[3][3] , \packet_addr[3][2] , 
        \packet_addr[3][1] , \packet_addr[3][0] }), .packet_addr_x_i({
        \packet_addr[3][7] , \packet_addr[3][6] , \packet_addr[3][5] , 
        \packet_addr[3][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[3]), 
        .east_req(\request[2][2] ), .local_req(\request[4][3] ) );
  dccl_5 dccl_l ( .packet_addr_y_i({\packet_addr[4][3] , \packet_addr[4][2] , 
        \packet_addr[4][1] , \packet_addr[4][0] }), .packet_addr_x_i({
        \packet_addr[4][7] , \packet_addr[4][6] , \packet_addr[4][5] , 
        \packet_addr[4][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[4]), 
        .north_req(\request[0][1] ), .east_req(\request[2][3] ), .south_req(
        \request[1][1] ), .west_req(\request[3][3] ) );
endmodule


module mux2_1_3 ( data0, data1, select0, select1, data_o );
  input [15:0] data0;
  input [15:0] data1;
  output [15:0] data_o;
  input select0, select1;
  wire   n1, n4, n5;

  AO22X1 U4 ( .IN1(data1[9]), .IN2(n5), .IN3(data0[9]), .IN4(n4), .Q(data_o[9]) );
  AO22X1 U5 ( .IN1(data1[8]), .IN2(n5), .IN3(data0[8]), .IN4(n4), .Q(data_o[8]) );
  AO22X1 U6 ( .IN1(data1[7]), .IN2(n5), .IN3(data0[7]), .IN4(n4), .Q(data_o[7]) );
  AO22X1 U7 ( .IN1(data1[6]), .IN2(n5), .IN3(data0[6]), .IN4(n4), .Q(data_o[6]) );
  AO22X1 U8 ( .IN1(data1[5]), .IN2(n5), .IN3(data0[5]), .IN4(n4), .Q(data_o[5]) );
  AO22X1 U9 ( .IN1(data1[4]), .IN2(n5), .IN3(data0[4]), .IN4(n4), .Q(data_o[4]) );
  AO22X1 U10 ( .IN1(data1[3]), .IN2(n5), .IN3(data0[3]), .IN4(n4), .Q(
        data_o[3]) );
  AO22X1 U11 ( .IN1(data1[2]), .IN2(n5), .IN3(data0[2]), .IN4(n4), .Q(
        data_o[2]) );
  AO22X1 U12 ( .IN1(data1[1]), .IN2(n5), .IN3(data0[1]), .IN4(n4), .Q(
        data_o[1]) );
  AO22X1 U13 ( .IN1(data1[15]), .IN2(n5), .IN3(data0[15]), .IN4(n4), .Q(
        data_o[15]) );
  AO22X1 U14 ( .IN1(data1[14]), .IN2(n5), .IN3(data0[14]), .IN4(n4), .Q(
        data_o[14]) );
  AO22X1 U15 ( .IN1(data1[13]), .IN2(n5), .IN3(data0[13]), .IN4(n4), .Q(
        data_o[13]) );
  AO22X1 U16 ( .IN1(data1[12]), .IN2(n5), .IN3(data0[12]), .IN4(n4), .Q(
        data_o[12]) );
  AO22X1 U17 ( .IN1(data1[11]), .IN2(n5), .IN3(data0[11]), .IN4(n4), .Q(
        data_o[11]) );
  AO22X1 U18 ( .IN1(data1[10]), .IN2(n5), .IN3(data0[10]), .IN4(n4), .Q(
        data_o[10]) );
  AO22X1 U19 ( .IN1(data1[0]), .IN2(n5), .IN3(data0[0]), .IN4(n4), .Q(
        data_o[0]) );
  INVX0 U2 ( .INP(select1), .ZN(n1) );
  AND2X1 U3 ( .IN1(select0), .IN2(n1), .Q(n4) );
  NOR2X0 U20 ( .IN1(n1), .IN2(select0), .QN(n5) );
endmodule


module mux2_1_2 ( data0, data1, select0, select1, data_o );
  input [15:0] data0;
  input [15:0] data1;
  output [15:0] data_o;
  input select0, select1;
  wire   n1, n4, n5;

  AO22X1 U4 ( .IN1(data1[9]), .IN2(n5), .IN3(data0[9]), .IN4(n4), .Q(data_o[9]) );
  AO22X1 U5 ( .IN1(data1[8]), .IN2(n5), .IN3(data0[8]), .IN4(n4), .Q(data_o[8]) );
  AO22X1 U6 ( .IN1(data1[7]), .IN2(n5), .IN3(data0[7]), .IN4(n4), .Q(data_o[7]) );
  AO22X1 U7 ( .IN1(data1[6]), .IN2(n5), .IN3(data0[6]), .IN4(n4), .Q(data_o[6]) );
  AO22X1 U8 ( .IN1(data1[5]), .IN2(n5), .IN3(data0[5]), .IN4(n4), .Q(data_o[5]) );
  AO22X1 U9 ( .IN1(data1[4]), .IN2(n5), .IN3(data0[4]), .IN4(n4), .Q(data_o[4]) );
  AO22X1 U10 ( .IN1(data1[3]), .IN2(n5), .IN3(data0[3]), .IN4(n4), .Q(
        data_o[3]) );
  AO22X1 U11 ( .IN1(data1[2]), .IN2(n5), .IN3(data0[2]), .IN4(n4), .Q(
        data_o[2]) );
  AO22X1 U12 ( .IN1(data1[1]), .IN2(n5), .IN3(data0[1]), .IN4(n4), .Q(
        data_o[1]) );
  AO22X1 U13 ( .IN1(data1[15]), .IN2(n5), .IN3(data0[15]), .IN4(n4), .Q(
        data_o[15]) );
  AO22X1 U14 ( .IN1(data1[14]), .IN2(n5), .IN3(data0[14]), .IN4(n4), .Q(
        data_o[14]) );
  AO22X1 U15 ( .IN1(data1[13]), .IN2(n5), .IN3(data0[13]), .IN4(n4), .Q(
        data_o[13]) );
  AO22X1 U16 ( .IN1(data1[12]), .IN2(n5), .IN3(data0[12]), .IN4(n4), .Q(
        data_o[12]) );
  AO22X1 U17 ( .IN1(data1[11]), .IN2(n5), .IN3(data0[11]), .IN4(n4), .Q(
        data_o[11]) );
  AO22X1 U18 ( .IN1(data1[10]), .IN2(n5), .IN3(data0[10]), .IN4(n4), .Q(
        data_o[10]) );
  AO22X1 U19 ( .IN1(data1[0]), .IN2(n5), .IN3(data0[0]), .IN4(n4), .Q(
        data_o[0]) );
  INVX0 U2 ( .INP(select1), .ZN(n1) );
  AND2X1 U3 ( .IN1(select0), .IN2(n1), .Q(n4) );
  NOR2X0 U20 ( .IN1(n1), .IN2(select0), .QN(n5) );
endmodule


module mux4_1_5 ( data0, data1, data2, data3, select0, select1, select2, 
        select3, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  input [15:0] data3;
  output [15:0] data_o;
  input select0, select1, select2, select3;
  wire   n1, n2, n3, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43;

  AO221X1 U5 ( .IN1(data1[9]), .IN2(n43), .IN3(data0[9]), .IN4(n42), .IN5(n41), 
        .Q(data_o[9]) );
  AO22X1 U6 ( .IN1(data2[9]), .IN2(n40), .IN3(data3[9]), .IN4(n39), .Q(n41) );
  AO221X1 U7 ( .IN1(data1[8]), .IN2(n43), .IN3(data0[8]), .IN4(n42), .IN5(n38), 
        .Q(data_o[8]) );
  AO22X1 U8 ( .IN1(data2[8]), .IN2(n40), .IN3(data3[8]), .IN4(n39), .Q(n38) );
  AO221X1 U9 ( .IN1(data1[7]), .IN2(n43), .IN3(data0[7]), .IN4(n42), .IN5(n37), 
        .Q(data_o[7]) );
  AO22X1 U10 ( .IN1(data2[7]), .IN2(n40), .IN3(data3[7]), .IN4(n39), .Q(n37)
         );
  AO221X1 U11 ( .IN1(data1[6]), .IN2(n43), .IN3(data0[6]), .IN4(n42), .IN5(n36), .Q(data_o[6]) );
  AO22X1 U12 ( .IN1(data2[6]), .IN2(n40), .IN3(data3[6]), .IN4(n39), .Q(n36)
         );
  AO221X1 U13 ( .IN1(data1[5]), .IN2(n43), .IN3(data0[5]), .IN4(n42), .IN5(n35), .Q(data_o[5]) );
  AO22X1 U14 ( .IN1(data2[5]), .IN2(n40), .IN3(data3[5]), .IN4(n39), .Q(n35)
         );
  AO221X1 U15 ( .IN1(data1[4]), .IN2(n43), .IN3(data0[4]), .IN4(n42), .IN5(n34), .Q(data_o[4]) );
  AO22X1 U16 ( .IN1(data2[4]), .IN2(n40), .IN3(data3[4]), .IN4(n39), .Q(n34)
         );
  AO221X1 U17 ( .IN1(data1[3]), .IN2(n43), .IN3(data0[3]), .IN4(n42), .IN5(n33), .Q(data_o[3]) );
  AO22X1 U18 ( .IN1(data2[3]), .IN2(n40), .IN3(data3[3]), .IN4(n39), .Q(n33)
         );
  AO221X1 U19 ( .IN1(data1[2]), .IN2(n43), .IN3(data0[2]), .IN4(n42), .IN5(n32), .Q(data_o[2]) );
  AO22X1 U20 ( .IN1(data2[2]), .IN2(n40), .IN3(data3[2]), .IN4(n39), .Q(n32)
         );
  AO221X1 U21 ( .IN1(data1[1]), .IN2(n43), .IN3(data0[1]), .IN4(n42), .IN5(n31), .Q(data_o[1]) );
  AO22X1 U22 ( .IN1(data2[1]), .IN2(n40), .IN3(data3[1]), .IN4(n39), .Q(n31)
         );
  AO221X1 U23 ( .IN1(data1[15]), .IN2(n43), .IN3(data0[15]), .IN4(n42), .IN5(
        n30), .Q(data_o[15]) );
  AO22X1 U24 ( .IN1(data2[15]), .IN2(n40), .IN3(data3[15]), .IN4(n39), .Q(n30)
         );
  AO221X1 U25 ( .IN1(data1[14]), .IN2(n43), .IN3(data0[14]), .IN4(n42), .IN5(
        n29), .Q(data_o[14]) );
  AO22X1 U26 ( .IN1(data2[14]), .IN2(n40), .IN3(data3[14]), .IN4(n39), .Q(n29)
         );
  AO221X1 U27 ( .IN1(data1[13]), .IN2(n43), .IN3(data0[13]), .IN4(n42), .IN5(
        n28), .Q(data_o[13]) );
  AO22X1 U28 ( .IN1(data2[13]), .IN2(n40), .IN3(data3[13]), .IN4(n39), .Q(n28)
         );
  AO221X1 U29 ( .IN1(data1[12]), .IN2(n43), .IN3(data0[12]), .IN4(n42), .IN5(
        n27), .Q(data_o[12]) );
  AO22X1 U30 ( .IN1(data2[12]), .IN2(n40), .IN3(data3[12]), .IN4(n39), .Q(n27)
         );
  AO221X1 U31 ( .IN1(data1[11]), .IN2(n43), .IN3(data0[11]), .IN4(n42), .IN5(
        n26), .Q(data_o[11]) );
  AO22X1 U32 ( .IN1(data2[11]), .IN2(n40), .IN3(data3[11]), .IN4(n39), .Q(n26)
         );
  AO221X1 U33 ( .IN1(data1[10]), .IN2(n43), .IN3(data0[10]), .IN4(n42), .IN5(
        n25), .Q(data_o[10]) );
  AO22X1 U34 ( .IN1(data2[10]), .IN2(n40), .IN3(data3[10]), .IN4(n39), .Q(n25)
         );
  AO221X1 U35 ( .IN1(data1[0]), .IN2(n43), .IN3(data0[0]), .IN4(n42), .IN5(n24), .Q(data_o[0]) );
  AO22X1 U36 ( .IN1(data2[0]), .IN2(n40), .IN3(data3[0]), .IN4(n39), .Q(n24)
         );
  INVX0 U2 ( .INP(select2), .ZN(n1) );
  NOR4X0 U3 ( .IN1(n1), .IN2(select0), .IN3(select1), .IN4(select3), .QN(n40)
         );
  AND4X1 U4 ( .IN1(select3), .IN2(n3), .IN3(n2), .IN4(n1), .Q(n39) );
  INVX0 U37 ( .INP(select0), .ZN(n3) );
  INVX0 U38 ( .INP(select1), .ZN(n2) );
  NOR4X0 U39 ( .IN1(n3), .IN2(select1), .IN3(select2), .IN4(select3), .QN(n42)
         );
  NOR4X0 U40 ( .IN1(n2), .IN2(select0), .IN3(select2), .IN4(select3), .QN(n43)
         );
endmodule


module mux4_1_4 ( data0, data1, data2, data3, select0, select1, select2, 
        select3, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  input [15:0] data3;
  output [15:0] data_o;
  input select0, select1, select2, select3;
  wire   n1, n2, n3, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43;

  AO221X1 U5 ( .IN1(data1[9]), .IN2(n43), .IN3(data0[9]), .IN4(n42), .IN5(n41), 
        .Q(data_o[9]) );
  AO22X1 U6 ( .IN1(data2[9]), .IN2(n40), .IN3(data3[9]), .IN4(n39), .Q(n41) );
  AO221X1 U7 ( .IN1(data1[8]), .IN2(n43), .IN3(data0[8]), .IN4(n42), .IN5(n38), 
        .Q(data_o[8]) );
  AO22X1 U8 ( .IN1(data2[8]), .IN2(n40), .IN3(data3[8]), .IN4(n39), .Q(n38) );
  AO221X1 U9 ( .IN1(data1[7]), .IN2(n43), .IN3(data0[7]), .IN4(n42), .IN5(n37), 
        .Q(data_o[7]) );
  AO22X1 U10 ( .IN1(data2[7]), .IN2(n40), .IN3(data3[7]), .IN4(n39), .Q(n37)
         );
  AO221X1 U11 ( .IN1(data1[6]), .IN2(n43), .IN3(data0[6]), .IN4(n42), .IN5(n36), .Q(data_o[6]) );
  AO22X1 U12 ( .IN1(data2[6]), .IN2(n40), .IN3(data3[6]), .IN4(n39), .Q(n36)
         );
  AO221X1 U13 ( .IN1(data1[5]), .IN2(n43), .IN3(data0[5]), .IN4(n42), .IN5(n35), .Q(data_o[5]) );
  AO22X1 U14 ( .IN1(data2[5]), .IN2(n40), .IN3(data3[5]), .IN4(n39), .Q(n35)
         );
  AO221X1 U15 ( .IN1(data1[4]), .IN2(n43), .IN3(data0[4]), .IN4(n42), .IN5(n34), .Q(data_o[4]) );
  AO22X1 U16 ( .IN1(data2[4]), .IN2(n40), .IN3(data3[4]), .IN4(n39), .Q(n34)
         );
  AO221X1 U17 ( .IN1(data1[3]), .IN2(n43), .IN3(data0[3]), .IN4(n42), .IN5(n33), .Q(data_o[3]) );
  AO22X1 U18 ( .IN1(data2[3]), .IN2(n40), .IN3(data3[3]), .IN4(n39), .Q(n33)
         );
  AO221X1 U19 ( .IN1(data1[2]), .IN2(n43), .IN3(data0[2]), .IN4(n42), .IN5(n32), .Q(data_o[2]) );
  AO22X1 U20 ( .IN1(data2[2]), .IN2(n40), .IN3(data3[2]), .IN4(n39), .Q(n32)
         );
  AO221X1 U21 ( .IN1(data1[1]), .IN2(n43), .IN3(data0[1]), .IN4(n42), .IN5(n31), .Q(data_o[1]) );
  AO22X1 U22 ( .IN1(data2[1]), .IN2(n40), .IN3(data3[1]), .IN4(n39), .Q(n31)
         );
  AO221X1 U23 ( .IN1(data1[15]), .IN2(n43), .IN3(data0[15]), .IN4(n42), .IN5(
        n30), .Q(data_o[15]) );
  AO22X1 U24 ( .IN1(data2[15]), .IN2(n40), .IN3(data3[15]), .IN4(n39), .Q(n30)
         );
  AO221X1 U25 ( .IN1(data1[14]), .IN2(n43), .IN3(data0[14]), .IN4(n42), .IN5(
        n29), .Q(data_o[14]) );
  AO22X1 U26 ( .IN1(data2[14]), .IN2(n40), .IN3(data3[14]), .IN4(n39), .Q(n29)
         );
  AO221X1 U27 ( .IN1(data1[13]), .IN2(n43), .IN3(data0[13]), .IN4(n42), .IN5(
        n28), .Q(data_o[13]) );
  AO22X1 U28 ( .IN1(data2[13]), .IN2(n40), .IN3(data3[13]), .IN4(n39), .Q(n28)
         );
  AO221X1 U29 ( .IN1(data1[12]), .IN2(n43), .IN3(data0[12]), .IN4(n42), .IN5(
        n27), .Q(data_o[12]) );
  AO22X1 U30 ( .IN1(data2[12]), .IN2(n40), .IN3(data3[12]), .IN4(n39), .Q(n27)
         );
  AO221X1 U31 ( .IN1(data1[11]), .IN2(n43), .IN3(data0[11]), .IN4(n42), .IN5(
        n26), .Q(data_o[11]) );
  AO22X1 U32 ( .IN1(data2[11]), .IN2(n40), .IN3(data3[11]), .IN4(n39), .Q(n26)
         );
  AO221X1 U33 ( .IN1(data1[10]), .IN2(n43), .IN3(data0[10]), .IN4(n42), .IN5(
        n25), .Q(data_o[10]) );
  AO22X1 U34 ( .IN1(data2[10]), .IN2(n40), .IN3(data3[10]), .IN4(n39), .Q(n25)
         );
  AO221X1 U35 ( .IN1(data1[0]), .IN2(n43), .IN3(data0[0]), .IN4(n42), .IN5(n24), .Q(data_o[0]) );
  AO22X1 U36 ( .IN1(data2[0]), .IN2(n40), .IN3(data3[0]), .IN4(n39), .Q(n24)
         );
  INVX0 U2 ( .INP(select2), .ZN(n1) );
  NOR4X0 U3 ( .IN1(n1), .IN2(select0), .IN3(select1), .IN4(select3), .QN(n40)
         );
  AND4X1 U4 ( .IN1(select3), .IN2(n3), .IN3(n2), .IN4(n1), .Q(n39) );
  INVX0 U37 ( .INP(select0), .ZN(n3) );
  INVX0 U38 ( .INP(select1), .ZN(n2) );
  NOR4X0 U39 ( .IN1(n3), .IN2(select1), .IN3(select2), .IN4(select3), .QN(n42)
         );
  NOR4X0 U40 ( .IN1(n2), .IN2(select0), .IN3(select2), .IN4(select3), .QN(n43)
         );
endmodule


module mux4_1_3 ( data0, data1, data2, data3, select0, select1, select2, 
        select3, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  input [15:0] data3;
  output [15:0] data_o;
  input select0, select1, select2, select3;
  wire   n1, n2, n3, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43;

  AO221X1 U5 ( .IN1(data1[9]), .IN2(n43), .IN3(data0[9]), .IN4(n42), .IN5(n41), 
        .Q(data_o[9]) );
  AO22X1 U6 ( .IN1(data2[9]), .IN2(n40), .IN3(data3[9]), .IN4(n39), .Q(n41) );
  AO221X1 U7 ( .IN1(data1[8]), .IN2(n43), .IN3(data0[8]), .IN4(n42), .IN5(n38), 
        .Q(data_o[8]) );
  AO22X1 U8 ( .IN1(data2[8]), .IN2(n40), .IN3(data3[8]), .IN4(n39), .Q(n38) );
  AO221X1 U9 ( .IN1(data1[7]), .IN2(n43), .IN3(data0[7]), .IN4(n42), .IN5(n37), 
        .Q(data_o[7]) );
  AO22X1 U10 ( .IN1(data2[7]), .IN2(n40), .IN3(data3[7]), .IN4(n39), .Q(n37)
         );
  AO221X1 U11 ( .IN1(data1[6]), .IN2(n43), .IN3(data0[6]), .IN4(n42), .IN5(n36), .Q(data_o[6]) );
  AO22X1 U12 ( .IN1(data2[6]), .IN2(n40), .IN3(data3[6]), .IN4(n39), .Q(n36)
         );
  AO221X1 U13 ( .IN1(data1[5]), .IN2(n43), .IN3(data0[5]), .IN4(n42), .IN5(n35), .Q(data_o[5]) );
  AO22X1 U14 ( .IN1(data2[5]), .IN2(n40), .IN3(data3[5]), .IN4(n39), .Q(n35)
         );
  AO221X1 U15 ( .IN1(data1[4]), .IN2(n43), .IN3(data0[4]), .IN4(n42), .IN5(n34), .Q(data_o[4]) );
  AO22X1 U16 ( .IN1(data2[4]), .IN2(n40), .IN3(data3[4]), .IN4(n39), .Q(n34)
         );
  AO221X1 U17 ( .IN1(data1[3]), .IN2(n43), .IN3(data0[3]), .IN4(n42), .IN5(n33), .Q(data_o[3]) );
  AO22X1 U18 ( .IN1(data2[3]), .IN2(n40), .IN3(data3[3]), .IN4(n39), .Q(n33)
         );
  AO221X1 U19 ( .IN1(data1[2]), .IN2(n43), .IN3(data0[2]), .IN4(n42), .IN5(n32), .Q(data_o[2]) );
  AO22X1 U20 ( .IN1(data2[2]), .IN2(n40), .IN3(data3[2]), .IN4(n39), .Q(n32)
         );
  AO221X1 U21 ( .IN1(data1[1]), .IN2(n43), .IN3(data0[1]), .IN4(n42), .IN5(n31), .Q(data_o[1]) );
  AO22X1 U22 ( .IN1(data2[1]), .IN2(n40), .IN3(data3[1]), .IN4(n39), .Q(n31)
         );
  AO221X1 U23 ( .IN1(data1[15]), .IN2(n43), .IN3(data0[15]), .IN4(n42), .IN5(
        n30), .Q(data_o[15]) );
  AO22X1 U24 ( .IN1(data2[15]), .IN2(n40), .IN3(data3[15]), .IN4(n39), .Q(n30)
         );
  AO221X1 U25 ( .IN1(data1[14]), .IN2(n43), .IN3(data0[14]), .IN4(n42), .IN5(
        n29), .Q(data_o[14]) );
  AO22X1 U26 ( .IN1(data2[14]), .IN2(n40), .IN3(data3[14]), .IN4(n39), .Q(n29)
         );
  AO221X1 U27 ( .IN1(data1[13]), .IN2(n43), .IN3(data0[13]), .IN4(n42), .IN5(
        n28), .Q(data_o[13]) );
  AO22X1 U28 ( .IN1(data2[13]), .IN2(n40), .IN3(data3[13]), .IN4(n39), .Q(n28)
         );
  AO221X1 U29 ( .IN1(data1[12]), .IN2(n43), .IN3(data0[12]), .IN4(n42), .IN5(
        n27), .Q(data_o[12]) );
  AO22X1 U30 ( .IN1(data2[12]), .IN2(n40), .IN3(data3[12]), .IN4(n39), .Q(n27)
         );
  AO221X1 U31 ( .IN1(data1[11]), .IN2(n43), .IN3(data0[11]), .IN4(n42), .IN5(
        n26), .Q(data_o[11]) );
  AO22X1 U32 ( .IN1(data2[11]), .IN2(n40), .IN3(data3[11]), .IN4(n39), .Q(n26)
         );
  AO221X1 U33 ( .IN1(data1[10]), .IN2(n43), .IN3(data0[10]), .IN4(n42), .IN5(
        n25), .Q(data_o[10]) );
  AO22X1 U34 ( .IN1(data2[10]), .IN2(n40), .IN3(data3[10]), .IN4(n39), .Q(n25)
         );
  AO221X1 U35 ( .IN1(data1[0]), .IN2(n43), .IN3(data0[0]), .IN4(n42), .IN5(n24), .Q(data_o[0]) );
  AO22X1 U36 ( .IN1(data2[0]), .IN2(n40), .IN3(data3[0]), .IN4(n39), .Q(n24)
         );
  INVX0 U2 ( .INP(select2), .ZN(n1) );
  NOR4X0 U3 ( .IN1(n1), .IN2(select0), .IN3(select1), .IN4(select3), .QN(n40)
         );
  AND4X1 U4 ( .IN1(select3), .IN2(n3), .IN3(n2), .IN4(n1), .Q(n39) );
  INVX0 U37 ( .INP(select0), .ZN(n3) );
  INVX0 U38 ( .INP(select1), .ZN(n2) );
  NOR4X0 U39 ( .IN1(n3), .IN2(select1), .IN3(select2), .IN4(select3), .QN(n42)
         );
  NOR4X0 U40 ( .IN1(n2), .IN2(select0), .IN3(select2), .IN4(select3), .QN(n43)
         );
endmodule



    module node5_NODE_X2_NODE_Y1I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__I_node_2_node_interface__I_node_3_node_interface__ ( 
        \clk.clk , \reset.reset , \local_node.clk , 
        \local_node.buffer_full_in , \local_node.buffer_full_out , 
        \local_node.receiving_data , \local_node.sending_data , 
        \local_node.data_in , \local_node.data_out , \node_0.clk , 
        \node_0.buffer_full_in , \node_0.buffer_full_out , 
        \node_0.receiving_data , \node_0.sending_data , \node_0.data_in , 
        \node_0.data_out , \node_1.clk , \node_1.buffer_full_in , 
        \node_1.buffer_full_out , \node_1.receiving_data , 
        \node_1.sending_data , \node_1.data_in , \node_1.data_out , 
        \node_2.clk , \node_2.buffer_full_in , \node_2.buffer_full_out , 
        \node_2.receiving_data , \node_2.sending_data , \node_2.data_in , 
        \node_2.data_out , \node_3.clk , \node_3.buffer_full_in , 
        \node_3.buffer_full_out , \node_3.receiving_data , 
        \node_3.sending_data , \node_3.data_in , \node_3.data_out  );
  input [15:0] \local_node.data_in ;
  output [15:0] \local_node.data_out ;
  input [15:0] \node_0.data_in ;
  output [15:0] \node_0.data_out ;
  input [15:0] \node_1.data_in ;
  output [15:0] \node_1.data_out ;
  input [15:0] \node_2.data_in ;
  output [15:0] \node_2.data_out ;
  input [15:0] \node_3.data_in ;
  output [15:0] \node_3.data_out ;
  input \clk.clk , \reset.reset , \local_node.buffer_full_in ,
         \local_node.receiving_data , \node_0.buffer_full_in ,
         \node_0.receiving_data , \node_1.buffer_full_in ,
         \node_1.receiving_data , \node_2.buffer_full_in ,
         \node_2.receiving_data , \node_3.buffer_full_in ,
         \node_3.receiving_data ;
  output \local_node.buffer_full_out , \local_node.sending_data ,
         \node_0.buffer_full_out , \node_0.sending_data ,
         \node_1.buffer_full_out , \node_1.sending_data ,
         \node_2.buffer_full_out , \node_2.sending_data ,
         \node_3.buffer_full_out , \node_3.sending_data ;
  inout \local_node.clk ,  \node_0.clk ,  \node_1.clk ,  \node_2.clk , 
     \node_3.clk ;
  wire   \buffer_out[4][15] , \buffer_out[4][14] , \buffer_out[4][13] ,
         \buffer_out[4][12] , \buffer_out[4][11] , \buffer_out[4][10] ,
         \buffer_out[4][9] , \buffer_out[4][8] , \buffer_out[4][7] ,
         \buffer_out[4][6] , \buffer_out[4][5] , \buffer_out[4][4] ,
         \buffer_out[4][3] , \buffer_out[4][2] , \buffer_out[4][1] ,
         \buffer_out[4][0] , \buffer_out[3][15] , \buffer_out[3][14] ,
         \buffer_out[3][13] , \buffer_out[3][12] , \buffer_out[3][11] ,
         \buffer_out[3][10] , \buffer_out[3][9] , \buffer_out[3][8] ,
         \buffer_out[3][7] , \buffer_out[3][6] , \buffer_out[3][5] ,
         \buffer_out[3][4] , \buffer_out[3][3] , \buffer_out[3][2] ,
         \buffer_out[3][1] , \buffer_out[3][0] , \buffer_out[2][15] ,
         \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] ,
         \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] ,
         \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] ,
         \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] ,
         \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] ,
         \buffer_out[1][15] , \buffer_out[1][14] , \buffer_out[1][13] ,
         \buffer_out[1][12] , \buffer_out[1][11] , \buffer_out[1][10] ,
         \buffer_out[1][9] , \buffer_out[1][8] , \buffer_out[1][7] ,
         \buffer_out[1][6] , \buffer_out[1][5] , \buffer_out[1][4] ,
         \buffer_out[1][3] , \buffer_out[1][2] , \buffer_out[1][1] ,
         \buffer_out[1][0] , \buffer_out[0][15] , \buffer_out[0][14] ,
         \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] ,
         \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] ,
         \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] ,
         \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] ,
         \buffer_out[0][1] , \buffer_out[0][0] , \next_buffer_out[4][15] ,
         \next_buffer_out[4][14] , \next_buffer_out[4][13] ,
         \next_buffer_out[4][12] , \next_buffer_out[4][11] ,
         \next_buffer_out[4][10] , \next_buffer_out[4][9] ,
         \next_buffer_out[4][8] , \next_buffer_out[4][7] ,
         \next_buffer_out[4][6] , \next_buffer_out[4][5] ,
         \next_buffer_out[4][4] , \next_buffer_out[4][3] ,
         \next_buffer_out[4][2] , \next_buffer_out[4][1] ,
         \next_buffer_out[4][0] , \next_buffer_out[3][15] ,
         \next_buffer_out[3][14] , \next_buffer_out[3][13] ,
         \next_buffer_out[3][12] , \next_buffer_out[3][11] ,
         \next_buffer_out[3][10] , \next_buffer_out[3][9] ,
         \next_buffer_out[3][8] , \next_buffer_out[3][7] ,
         \next_buffer_out[3][6] , \next_buffer_out[3][5] ,
         \next_buffer_out[3][4] , \next_buffer_out[3][3] ,
         \next_buffer_out[3][2] , \next_buffer_out[3][1] ,
         \next_buffer_out[3][0] , \next_buffer_out[2][15] ,
         \next_buffer_out[2][14] , \next_buffer_out[2][13] ,
         \next_buffer_out[2][12] , \next_buffer_out[2][11] ,
         \next_buffer_out[2][10] , \next_buffer_out[2][9] ,
         \next_buffer_out[2][8] , \next_buffer_out[2][7] ,
         \next_buffer_out[2][6] , \next_buffer_out[2][5] ,
         \next_buffer_out[2][4] , \next_buffer_out[2][3] ,
         \next_buffer_out[2][2] , \next_buffer_out[2][1] ,
         \next_buffer_out[2][0] , \next_buffer_out[1][15] ,
         \next_buffer_out[1][14] , \next_buffer_out[1][13] ,
         \next_buffer_out[1][12] , \next_buffer_out[1][11] ,
         \next_buffer_out[1][10] , \next_buffer_out[1][9] ,
         \next_buffer_out[1][8] , \next_buffer_out[1][7] ,
         \next_buffer_out[1][6] , \next_buffer_out[1][5] ,
         \next_buffer_out[1][4] , \next_buffer_out[1][3] ,
         \next_buffer_out[1][2] , \next_buffer_out[1][1] ,
         \next_buffer_out[1][0] , \next_buffer_out[0][15] ,
         \next_buffer_out[0][14] , \next_buffer_out[0][13] ,
         \next_buffer_out[0][12] , \next_buffer_out[0][11] ,
         \next_buffer_out[0][10] , \next_buffer_out[0][9] ,
         \next_buffer_out[0][8] , \next_buffer_out[0][7] ,
         \next_buffer_out[0][6] , \next_buffer_out[0][5] ,
         \next_buffer_out[0][4] , \next_buffer_out[0][3] ,
         \next_buffer_out[0][2] , \next_buffer_out[0][1] ,
         \next_buffer_out[0][0] ;
  wire   [4:0] buffer_full_in;
  wire   [4:0] receiving_data;
  wire   [4:0] pop_v;
  wire   [4:0] data_valid;
  wire   [4:0] next_data_valid;
  wire   [1:0] grant_0;
  wire   [1:0] grant_1;
  wire   [3:0] grant_2;
  wire   [3:0] grant_3;
  wire   [3:0] grant_4;
  tri   \local_node.buffer_full_in ;
  tri   \local_node.buffer_full_out ;
  tri   \local_node.receiving_data ;
  tri   \local_node.sending_data ;
  tri   [15:0] \local_node.data_in ;
  tri   [15:0] \local_node.data_out ;

  converter_in_I_n_node_interface_dut__3 c0 ( .\n.buffer_full_in (
        \node_0.buffer_full_in ), .\n.receiving_data (\node_0.receiving_data ), 
        .\n.data_in (\node_0.data_in ), .\n.buffer_full_out (
        \node_0.buffer_full_out ), .\n.sending_data (\node_0.sending_data ), 
        .\n.data_out (\node_0.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_out_I_n_node_interface_dut_ c1 ( .\n.buffer_full_in (
        \node_1.buffer_full_in ), .\n.receiving_data (\node_1.receiving_data ), 
        .\n.data_in (\node_1.data_in ), .\n.buffer_full_out (
        \node_1.buffer_full_out ), .\n.sending_data (\node_1.sending_data ), 
        .\n.data_out (\node_1.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_in_I_n_node_interface_dut__2 c2 ( .\n.buffer_full_in (
        \node_2.buffer_full_in ), .\n.receiving_data (\node_2.receiving_data ), 
        .\n.data_in (\node_2.data_in ), .\n.buffer_full_out (
        \node_2.buffer_full_out ), .\n.sending_data (\node_2.sending_data ), 
        .\n.data_out (\node_2.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_out_I_n_node_interface_dut_ c3 ( .\n.buffer_full_in (
        \node_3.buffer_full_in ), .\n.receiving_data (\node_3.receiving_data ), 
        .\n.data_in (\node_3.data_in ), .\n.buffer_full_out (
        \node_3.buffer_full_out ), .\n.sending_data (\node_3.sending_data ), 
        .\n.data_out (\node_3.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_out_I_n_node_interface_dut_ c4 ( .\n.buffer_full_in (
        \local_node.buffer_full_in ), .\n.receiving_data (
        \local_node.receiving_data ), .\n.data_in (\local_node.data_in ), 
        .\n.buffer_full_out (\local_node.buffer_full_out ), .\n.sending_data (
        \local_node.sending_data ), .\n.data_out (\local_node.data_out ), 
        .buffer_full_in(1'b0), .receiving_data(1'b0), .data_in({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  fifo_kev_9 \genblk1[0].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[0]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[0]), .data_out({\buffer_out[0][15] , 
        \buffer_out[0][14] , \buffer_out[0][13] , \buffer_out[0][12] , 
        \buffer_out[0][11] , \buffer_out[0][10] , \buffer_out[0][9] , 
        \buffer_out[0][8] , \buffer_out[0][7] , \buffer_out[0][6] , 
        \buffer_out[0][5] , \buffer_out[0][4] , \buffer_out[0][3] , 
        \buffer_out[0][2] , \buffer_out[0][1] , \buffer_out[0][0] }), 
        .next_data_out({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] , 
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .next_data_valid(
        next_data_valid[0]) );
  address_counter_9 \genblk1[0].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] }), 
        .buffer_data_valid(next_data_valid[0]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .buffer_pop(
        pop_v[0]), .receiving_data(1'b0) );
  fifo_kev_8 \genblk1[1].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[1]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[1]), .data_out({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), 
        .next_data_out({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] , 
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .next_data_valid(
        next_data_valid[1]) );
  address_counter_8 \genblk1[1].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] }), 
        .buffer_data_valid(next_data_valid[1]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .buffer_pop(
        pop_v[1]), .receiving_data(1'b0) );
  fifo_kev_7 \genblk1[2].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[2]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[2]), .data_out({\buffer_out[2][15] , 
        \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] , 
        \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] , 
        \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] , 
        \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] , 
        \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] }), 
        .next_data_out({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] , 
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .next_data_valid(
        next_data_valid[2]) );
  address_counter_7 \genblk1[2].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] }), 
        .buffer_data_valid(next_data_valid[2]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .buffer_pop(
        pop_v[2]), .receiving_data(1'b0) );
  fifo_kev_6 \genblk1[3].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[3]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[3]), .data_out({\buffer_out[3][15] , 
        \buffer_out[3][14] , \buffer_out[3][13] , \buffer_out[3][12] , 
        \buffer_out[3][11] , \buffer_out[3][10] , \buffer_out[3][9] , 
        \buffer_out[3][8] , \buffer_out[3][7] , \buffer_out[3][6] , 
        \buffer_out[3][5] , \buffer_out[3][4] , \buffer_out[3][3] , 
        \buffer_out[3][2] , \buffer_out[3][1] , \buffer_out[3][0] }), 
        .next_data_out({\next_buffer_out[3][15] , \next_buffer_out[3][14] , 
        \next_buffer_out[3][13] , \next_buffer_out[3][12] , 
        \next_buffer_out[3][11] , \next_buffer_out[3][10] , 
        \next_buffer_out[3][9] , \next_buffer_out[3][8] , 
        \next_buffer_out[3][7] , \next_buffer_out[3][6] , 
        \next_buffer_out[3][5] , \next_buffer_out[3][4] , 
        \next_buffer_out[3][3] , \next_buffer_out[3][2] , 
        \next_buffer_out[3][1] , \next_buffer_out[3][0] }), .next_data_valid(
        next_data_valid[3]) );
  address_counter_6 \genblk1[3].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[3][15] , \next_buffer_out[3][14] , 
        \next_buffer_out[3][13] , \next_buffer_out[3][12] , 
        \next_buffer_out[3][11] , \next_buffer_out[3][10] , 
        \next_buffer_out[3][9] , \next_buffer_out[3][8] }), 
        .buffer_data_valid(next_data_valid[3]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[3][7] , \next_buffer_out[3][6] , 
        \next_buffer_out[3][5] , \next_buffer_out[3][4] , 
        \next_buffer_out[3][3] , \next_buffer_out[3][2] , 
        \next_buffer_out[3][1] , \next_buffer_out[3][0] }), .buffer_pop(
        pop_v[3]), .receiving_data(1'b0) );
  fifo_kev_5 \genblk1[4].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[4]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[4]), .data_out({\buffer_out[4][15] , 
        \buffer_out[4][14] , \buffer_out[4][13] , \buffer_out[4][12] , 
        \buffer_out[4][11] , \buffer_out[4][10] , \buffer_out[4][9] , 
        \buffer_out[4][8] , \buffer_out[4][7] , \buffer_out[4][6] , 
        \buffer_out[4][5] , \buffer_out[4][4] , \buffer_out[4][3] , 
        \buffer_out[4][2] , \buffer_out[4][1] , \buffer_out[4][0] }), 
        .next_data_out({\next_buffer_out[4][15] , \next_buffer_out[4][14] , 
        \next_buffer_out[4][13] , \next_buffer_out[4][12] , 
        \next_buffer_out[4][11] , \next_buffer_out[4][10] , 
        \next_buffer_out[4][9] , \next_buffer_out[4][8] , 
        \next_buffer_out[4][7] , \next_buffer_out[4][6] , 
        \next_buffer_out[4][5] , \next_buffer_out[4][4] , 
        \next_buffer_out[4][3] , \next_buffer_out[4][2] , 
        \next_buffer_out[4][1] , \next_buffer_out[4][0] }), .next_data_valid(
        next_data_valid[4]) );
  address_counter_5 \genblk1[4].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[4][15] , \next_buffer_out[4][14] , 
        \next_buffer_out[4][13] , \next_buffer_out[4][12] , 
        \next_buffer_out[4][11] , \next_buffer_out[4][10] , 
        \next_buffer_out[4][9] , \next_buffer_out[4][8] }), 
        .buffer_data_valid(next_data_valid[4]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[4][7] , \next_buffer_out[4][6] , 
        \next_buffer_out[4][5] , \next_buffer_out[4][4] , 
        \next_buffer_out[4][3] , \next_buffer_out[4][2] , 
        \next_buffer_out[4][1] , \next_buffer_out[4][0] }), .buffer_pop(
        pop_v[4]), .receiving_data(1'b0) );
  controller5_1 ctrl5 ( .clk(\clk.clk ), .rst(\reset.reset ), .packet_addr({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .local_addr({1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b1}), .packet_valid(data_valid), .buffer_full_in({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .grant_0(grant_0), .grant_1(grant_1), 
        .grant_2(grant_2), .grant_3(grant_3), .grant_4(grant_4), .pop_v(pop_v)
         );
  mux2_1_3 mux_n ( .data0({\buffer_out[1][15] , \buffer_out[1][14] , 
        \buffer_out[1][13] , \buffer_out[1][12] , \buffer_out[1][11] , 
        \buffer_out[1][10] , \buffer_out[1][9] , \buffer_out[1][8] , 
        \buffer_out[1][7] , \buffer_out[1][6] , \buffer_out[1][5] , 
        \buffer_out[1][4] , \buffer_out[1][3] , \buffer_out[1][2] , 
        \buffer_out[1][1] , \buffer_out[1][0] }), .data1({\buffer_out[4][15] , 
        \buffer_out[4][14] , \buffer_out[4][13] , \buffer_out[4][12] , 
        \buffer_out[4][11] , \buffer_out[4][10] , \buffer_out[4][9] , 
        \buffer_out[4][8] , \buffer_out[4][7] , \buffer_out[4][6] , 
        \buffer_out[4][5] , \buffer_out[4][4] , \buffer_out[4][3] , 
        \buffer_out[4][2] , \buffer_out[4][1] , \buffer_out[4][0] }), 
        .select0(grant_0[0]), .select1(grant_0[1]) );
  mux2_1_2 mux_s ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[4][15] , 
        \buffer_out[4][14] , \buffer_out[4][13] , \buffer_out[4][12] , 
        \buffer_out[4][11] , \buffer_out[4][10] , \buffer_out[4][9] , 
        \buffer_out[4][8] , \buffer_out[4][7] , \buffer_out[4][6] , 
        \buffer_out[4][5] , \buffer_out[4][4] , \buffer_out[4][3] , 
        \buffer_out[4][2] , \buffer_out[4][1] , \buffer_out[4][0] }), 
        .select0(grant_1[0]), .select1(grant_1[1]) );
  mux4_1_5 mux_e ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[3][15] , \buffer_out[3][14] , \buffer_out[3][13] , 
        \buffer_out[3][12] , \buffer_out[3][11] , \buffer_out[3][10] , 
        \buffer_out[3][9] , \buffer_out[3][8] , \buffer_out[3][7] , 
        \buffer_out[3][6] , \buffer_out[3][5] , \buffer_out[3][4] , 
        \buffer_out[3][3] , \buffer_out[3][2] , \buffer_out[3][1] , 
        \buffer_out[3][0] }), .data3({\buffer_out[4][15] , \buffer_out[4][14] , 
        \buffer_out[4][13] , \buffer_out[4][12] , \buffer_out[4][11] , 
        \buffer_out[4][10] , \buffer_out[4][9] , \buffer_out[4][8] , 
        \buffer_out[4][7] , \buffer_out[4][6] , \buffer_out[4][5] , 
        \buffer_out[4][4] , \buffer_out[4][3] , \buffer_out[4][2] , 
        \buffer_out[4][1] , \buffer_out[4][0] }), .select0(grant_2[0]), 
        .select1(grant_2[1]), .select2(grant_2[2]), .select3(grant_2[3]) );
  mux4_1_4 mux_w ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[2][15] , \buffer_out[2][14] , \buffer_out[2][13] , 
        \buffer_out[2][12] , \buffer_out[2][11] , \buffer_out[2][10] , 
        \buffer_out[2][9] , \buffer_out[2][8] , \buffer_out[2][7] , 
        \buffer_out[2][6] , \buffer_out[2][5] , \buffer_out[2][4] , 
        \buffer_out[2][3] , \buffer_out[2][2] , \buffer_out[2][1] , 
        \buffer_out[2][0] }), .data3({\buffer_out[4][15] , \buffer_out[4][14] , 
        \buffer_out[4][13] , \buffer_out[4][12] , \buffer_out[4][11] , 
        \buffer_out[4][10] , \buffer_out[4][9] , \buffer_out[4][8] , 
        \buffer_out[4][7] , \buffer_out[4][6] , \buffer_out[4][5] , 
        \buffer_out[4][4] , \buffer_out[4][3] , \buffer_out[4][2] , 
        \buffer_out[4][1] , \buffer_out[4][0] }), .select0(grant_3[0]), 
        .select1(grant_3[1]), .select2(grant_3[2]), .select3(grant_3[3]) );
  mux4_1_3 mux_l ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[2][15] , \buffer_out[2][14] , \buffer_out[2][13] , 
        \buffer_out[2][12] , \buffer_out[2][11] , \buffer_out[2][10] , 
        \buffer_out[2][9] , \buffer_out[2][8] , \buffer_out[2][7] , 
        \buffer_out[2][6] , \buffer_out[2][5] , \buffer_out[2][4] , 
        \buffer_out[2][3] , \buffer_out[2][2] , \buffer_out[2][1] , 
        \buffer_out[2][0] }), .data3({\buffer_out[3][15] , \buffer_out[3][14] , 
        \buffer_out[3][13] , \buffer_out[3][12] , \buffer_out[3][11] , 
        \buffer_out[3][10] , \buffer_out[3][9] , \buffer_out[3][8] , 
        \buffer_out[3][7] , \buffer_out[3][6] , \buffer_out[3][5] , 
        \buffer_out[3][4] , \buffer_out[3][3] , \buffer_out[3][2] , 
        \buffer_out[3][1] , \buffer_out[3][0] }), .select0(grant_4[0]), 
        .select1(grant_4[1]), .select2(grant_4[2]), .select3(grant_4[3]) );
endmodule


module converter_in_I_n_node_interface_dut__1 ( \n.buffer_full_in , 
        \n.receiving_data , \n.data_in , \n.buffer_full_out , \n.sending_data , 
        \n.data_out , buffer_full_out, sending_data, data_out, buffer_full_in, 
        receiving_data, data_in );
  input [15:0] \n.data_in ;
  output [15:0] \n.data_out ;
  output [15:0] data_out;
  input [15:0] data_in;
  input \n.buffer_full_in , \n.receiving_data , buffer_full_in, receiving_data;
  output \n.buffer_full_out , \n.sending_data , buffer_full_out, sending_data;
  wire   \n.buffer_full_in , \n.receiving_data , buffer_full_in,
         receiving_data;
  assign buffer_full_out = \n.buffer_full_in ;
  assign sending_data = \n.receiving_data ;
  assign data_out[15] = \n.data_in  [15];
  assign data_out[14] = \n.data_in  [14];
  assign data_out[13] = \n.data_in  [13];
  assign data_out[12] = \n.data_in  [12];
  assign data_out[11] = \n.data_in  [11];
  assign data_out[10] = \n.data_in  [10];
  assign data_out[9] = \n.data_in  [9];
  assign data_out[8] = \n.data_in  [8];
  assign data_out[7] = \n.data_in  [7];
  assign data_out[6] = \n.data_in  [6];
  assign data_out[5] = \n.data_in  [5];
  assign data_out[4] = \n.data_in  [4];
  assign data_out[3] = \n.data_in  [3];
  assign data_out[2] = \n.data_in  [2];
  assign data_out[1] = \n.data_in  [1];
  assign data_out[0] = \n.data_in  [0];
  assign \n.buffer_full_out  = buffer_full_in;
  assign \n.sending_data  = receiving_data;
  assign \n.data_out  [15] = data_in[15];
  assign \n.data_out  [14] = data_in[14];
  assign \n.data_out  [13] = data_in[13];
  assign \n.data_out  [12] = data_in[12];
  assign \n.data_out  [11] = data_in[11];
  assign \n.data_out  [10] = data_in[10];
  assign \n.data_out  [9] = data_in[9];
  assign \n.data_out  [8] = data_in[8];
  assign \n.data_out  [7] = data_in[7];
  assign \n.data_out  [6] = data_in[6];
  assign \n.data_out  [5] = data_in[5];
  assign \n.data_out  [4] = data_in[4];
  assign \n.data_out  [3] = data_in[3];
  assign \n.data_out  [2] = data_in[2];
  assign \n.data_out  [1] = data_in[1];
  assign \n.data_out  [0] = data_in[0];

endmodule


module converter_in_I_n_node_interface_dut__0 ( \n.buffer_full_in , 
        \n.receiving_data , \n.data_in , \n.buffer_full_out , \n.sending_data , 
        \n.data_out , buffer_full_out, sending_data, data_out, buffer_full_in, 
        receiving_data, data_in );
  input [15:0] \n.data_in ;
  output [15:0] \n.data_out ;
  output [15:0] data_out;
  input [15:0] data_in;
  input \n.buffer_full_in , \n.receiving_data , buffer_full_in, receiving_data;
  output \n.buffer_full_out , \n.sending_data , buffer_full_out, sending_data;
  wire   \n.buffer_full_in , \n.receiving_data , buffer_full_in,
         receiving_data;
  assign buffer_full_out = \n.buffer_full_in ;
  assign sending_data = \n.receiving_data ;
  assign data_out[15] = \n.data_in  [15];
  assign data_out[14] = \n.data_in  [14];
  assign data_out[13] = \n.data_in  [13];
  assign data_out[12] = \n.data_in  [12];
  assign data_out[11] = \n.data_in  [11];
  assign data_out[10] = \n.data_in  [10];
  assign data_out[9] = \n.data_in  [9];
  assign data_out[8] = \n.data_in  [8];
  assign data_out[7] = \n.data_in  [7];
  assign data_out[6] = \n.data_in  [6];
  assign data_out[5] = \n.data_in  [5];
  assign data_out[4] = \n.data_in  [4];
  assign data_out[3] = \n.data_in  [3];
  assign data_out[2] = \n.data_in  [2];
  assign data_out[1] = \n.data_in  [1];
  assign data_out[0] = \n.data_in  [0];
  assign \n.buffer_full_out  = buffer_full_in;
  assign \n.sending_data  = receiving_data;
  assign \n.data_out  [15] = data_in[15];
  assign \n.data_out  [14] = data_in[14];
  assign \n.data_out  [13] = data_in[13];
  assign \n.data_out  [12] = data_in[12];
  assign \n.data_out  [11] = data_in[11];
  assign \n.data_out  [10] = data_in[10];
  assign \n.data_out  [9] = data_in[9];
  assign \n.data_out  [8] = data_in[8];
  assign \n.data_out  [7] = data_in[7];
  assign \n.data_out  [6] = data_in[6];
  assign \n.data_out  [5] = data_in[5];
  assign \n.data_out  [4] = data_in[4];
  assign \n.data_out  [3] = data_in[3];
  assign \n.data_out  [2] = data_in[2];
  assign \n.data_out  [1] = data_in[1];
  assign \n.data_out  [0] = data_in[0];

endmodule


module fifo_kev_4 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_9 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_4 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_9 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, n15, 
        n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_8 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_4 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_8 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, n15, 
        n13, n11, n9, n7, n5}) );
endmodule


module address_counter_4_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_4 ( clk, rst, interface_flit_length, buffer_flit_length, 
        buffer_data_valid, interface_flit_address, buffer_flit_address, 
        buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_4 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_4 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_4_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), .SUM(
        {SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_3 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_7 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_3 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_7 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, n15, 
        n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_6 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_3 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_6 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, n15, 
        n13, n11, n9, n7, n5}) );
endmodule


module address_counter_3_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_3 ( clk, rst, interface_flit_length, buffer_flit_length, 
        buffer_data_valid, interface_flit_address, buffer_flit_address, 
        buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_3 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_3 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_3_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), .SUM(
        {SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_2 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_5 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_2 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_5 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, n15, 
        n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_4 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_2 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_4 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, n15, 
        n13, n11, n9, n7, n5}) );
endmodule


module address_counter_2_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_2 ( clk, rst, interface_flit_length, buffer_flit_length, 
        buffer_data_valid, interface_flit_address, buffer_flit_address, 
        buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_2 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_2 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_2_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), .SUM(
        {SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_1 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_3 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_1 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_3 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, n15, 
        n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_2 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_1 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_2 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, n15, 
        n13, n11, n9, n7, n5}) );
endmodule


module address_counter_1_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_1 ( clk, rst, interface_flit_length, buffer_flit_length, 
        buffer_data_valid, interface_flit_address, buffer_flit_address, 
        buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_1 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_1 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_1_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), .SUM(
        {SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module fifo_kev_0 ( clk, rst, push_req, pop_req, data_in, full, data_valid, 
        data_out, next_data_out, next_data_valid );
  input [15:0] data_in;
  output [15:0] data_out;
  output [15:0] next_data_out;
  input clk, rst, push_req, pop_req;
  output full, data_valid, next_data_valid;
  wire   head_empty, fifo_empty, n1, n3, n4, n12, n13, n14, n15, n16, n17;
  wire   [15:0] head_wrdata;

  OR4X1 U10 ( .IN1(n17), .IN2(n12), .IN3(head_empty), .IN4(full), .Q(n14) );
  AO22X1 U11 ( .IN1(data_valid), .IN2(n4), .IN3(n16), .IN4(n12), .Q(n13) );
  AO22X1 U12 ( .IN1(data_in[9]), .IN2(n3), .IN3(next_data_out[9]), .IN4(n15), 
        .Q(head_wrdata[9]) );
  AO22X1 U13 ( .IN1(data_in[8]), .IN2(n3), .IN3(next_data_out[8]), .IN4(n15), 
        .Q(head_wrdata[8]) );
  AO22X1 U14 ( .IN1(data_in[7]), .IN2(n3), .IN3(next_data_out[7]), .IN4(n15), 
        .Q(head_wrdata[7]) );
  AO22X1 U15 ( .IN1(data_in[6]), .IN2(n3), .IN3(next_data_out[6]), .IN4(n15), 
        .Q(head_wrdata[6]) );
  AO22X1 U16 ( .IN1(data_in[5]), .IN2(n3), .IN3(next_data_out[5]), .IN4(n15), 
        .Q(head_wrdata[5]) );
  AO22X1 U17 ( .IN1(data_in[4]), .IN2(n3), .IN3(next_data_out[4]), .IN4(n15), 
        .Q(head_wrdata[4]) );
  AO22X1 U18 ( .IN1(data_in[3]), .IN2(n3), .IN3(next_data_out[3]), .IN4(n15), 
        .Q(head_wrdata[3]) );
  AO22X1 U19 ( .IN1(data_in[2]), .IN2(n3), .IN3(next_data_out[2]), .IN4(n15), 
        .Q(head_wrdata[2]) );
  AO22X1 U20 ( .IN1(data_in[1]), .IN2(n3), .IN3(next_data_out[1]), .IN4(n15), 
        .Q(head_wrdata[1]) );
  AO22X1 U21 ( .IN1(data_in[15]), .IN2(n3), .IN3(next_data_out[15]), .IN4(n15), 
        .Q(head_wrdata[15]) );
  AO22X1 U22 ( .IN1(data_in[14]), .IN2(n3), .IN3(next_data_out[14]), .IN4(n15), 
        .Q(head_wrdata[14]) );
  AO22X1 U23 ( .IN1(data_in[13]), .IN2(n3), .IN3(next_data_out[13]), .IN4(n15), 
        .Q(head_wrdata[13]) );
  AO22X1 U24 ( .IN1(data_in[12]), .IN2(n3), .IN3(next_data_out[12]), .IN4(n15), 
        .Q(head_wrdata[12]) );
  AO22X1 U25 ( .IN1(data_in[11]), .IN2(n3), .IN3(next_data_out[11]), .IN4(n15), 
        .Q(head_wrdata[11]) );
  AO22X1 U26 ( .IN1(data_in[10]), .IN2(n3), .IN3(next_data_out[10]), .IN4(n15), 
        .Q(head_wrdata[10]) );
  AO22X1 U27 ( .IN1(data_in[0]), .IN2(n3), .IN3(next_data_out[0]), .IN4(n15), 
        .Q(head_wrdata[0]) );
  OA22X1 U2 ( .IN1(n12), .IN2(data_valid), .IN3(n4), .IN4(next_data_valid), 
        .Q(n15) );
  INVX0 U3 ( .INP(n15), .ZN(n3) );
  INVX0 U4 ( .INP(fifo_empty), .ZN(next_data_valid) );
  INVX0 U5 ( .INP(head_empty), .ZN(data_valid) );
  INVX0 U6 ( .INP(push_req), .ZN(n12) );
  NOR2X0 U7 ( .IN1(next_data_valid), .IN2(n4), .QN(n17) );
  INVX0 U8 ( .INP(pop_req), .ZN(n4) );
  NAND2X1 U9 ( .IN1(pop_req), .IN2(next_data_valid), .QN(n16) );
  INVX0 U28 ( .INP(rst), .ZN(n1) );
  DW_fifo_s1_sf_width16_depth2_ae_level1_af_level1_err_mode1_rst_mode1 buffer_head ( 
        .clk(clk), .rst_n(n1), .push_req_n(n13), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(head_wrdata), .empty(head_empty), .peek_out(data_out) );
  DW_fifo_s1_sf_width16_depth4_ae_level1_af_level1_err_mode1_rst_mode1 buffer ( 
        .clk(clk), .rst_n(n1), .push_req_n(n14), .pop_req_n(n4), .diag_n(1'b1), 
        .data_in(data_in), .empty(fifo_empty), .full(full), .peek_out(
        next_data_out) );
endmodule


module flipflop_BITS8_1 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS8_0 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_1 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, n15, 
        n13, n11, n9, n7, n5}) );
endmodule


module flipflop_BITS8_0 ( clk, data_i, data_o );
  input [7:0] data_i;
  output [7:0] data_o;
  input clk;


  DFFX1 \data_o_reg[7]  ( .D(data_i[7]), .CLK(clk), .Q(data_o[7]) );
  DFFX1 \data_o_reg[6]  ( .D(data_i[6]), .CLK(clk), .Q(data_o[6]) );
  DFFX1 \data_o_reg[5]  ( .D(data_i[5]), .CLK(clk), .Q(data_o[5]) );
  DFFX1 \data_o_reg[4]  ( .D(data_i[4]), .CLK(clk), .Q(data_o[4]) );
  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_8_0 ( clk, enable_i, reset, data_i, data_o );
  input [7:0] data_i;
  input [7:0] data_o;
  input clk, enable_i, reset;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n1, n5, n7, n9, n11, n13, n15,
         n17, n19, n20, n21;
  wire   [7:0] write_data;

  AO22X1 U5 ( .IN1(data_i[7]), .IN2(n21), .IN3(n22), .IN4(n20), .Q(
        write_data[7]) );
  AO22X1 U6 ( .IN1(data_i[6]), .IN2(n21), .IN3(n23), .IN4(n20), .Q(
        write_data[6]) );
  AO22X1 U7 ( .IN1(data_i[5]), .IN2(n21), .IN3(n24), .IN4(n20), .Q(
        write_data[5]) );
  AO22X1 U8 ( .IN1(data_i[4]), .IN2(n21), .IN3(n25), .IN4(n20), .Q(
        write_data[4]) );
  AO22X1 U9 ( .IN1(data_i[3]), .IN2(n21), .IN3(n26), .IN4(n20), .Q(
        write_data[3]) );
  AO22X1 U10 ( .IN1(data_i[2]), .IN2(n21), .IN3(n27), .IN4(n20), .Q(
        write_data[2]) );
  AO22X1 U11 ( .IN1(data_i[1]), .IN2(n21), .IN3(n28), .IN4(n20), .Q(
        write_data[1]) );
  AO22X1 U12 ( .IN1(data_i[0]), .IN2(n21), .IN3(n29), .IN4(n20), .Q(
        write_data[0]) );
  NOR2X0 U2 ( .IN1(n1), .IN2(reset), .QN(n21) );
  INVX0 U3 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U4 ( .IN1(enable_i), .IN2(reset), .QN(n20) );
  AND2X1 U13 ( .IN1(data_o[7]), .IN2(n19), .Q(n22) );
  AND2X1 U14 ( .IN1(data_o[6]), .IN2(n17), .Q(n23) );
  AND2X1 U15 ( .IN1(data_o[5]), .IN2(n15), .Q(n24) );
  AND2X1 U16 ( .IN1(data_o[4]), .IN2(n13), .Q(n25) );
  AND2X1 U17 ( .IN1(data_o[3]), .IN2(n11), .Q(n26) );
  AND2X1 U18 ( .IN1(data_o[2]), .IN2(n9), .Q(n27) );
  AND2X1 U19 ( .IN1(data_o[1]), .IN2(n7), .Q(n28) );
  AND2X1 U20 ( .IN1(data_o[0]), .IN2(n5), .Q(n29) );
  flipflop_BITS8_0 FF ( .clk(clk), .data_i(write_data), .data_o({n19, n17, n15, 
        n13, n11, n9, n7, n5}) );
endmodule


module address_counter_0_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module address_counter_0 ( clk, rst, interface_flit_length, buffer_flit_length, 
        buffer_data_valid, interface_flit_address, buffer_flit_address, 
        buffer_pop, receiving_data, flit_address_o );
  input [7:0] interface_flit_length;
  input [7:0] buffer_flit_length;
  input [7:0] interface_flit_address;
  input [7:0] buffer_flit_address;
  output [7:0] flit_address_o;
  input clk, rst, buffer_data_valid, buffer_pop, receiving_data;
  wire   is_address, N12, N13, N14, N15, N16, N17, N18, N19, n1;
  wire   [7:0] current_count;
  wire   [7:0] next_count;
  wire   [7:0] flit_address;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign flit_address_o[0] = 1'b0;
  assign flit_address_o[1] = 1'b0;
  assign flit_address_o[2] = 1'b0;
  assign flit_address_o[3] = 1'b0;
  assign flit_address_o[4] = 1'b0;
  assign flit_address_o[5] = 1'b0;
  assign flit_address_o[6] = 1'b0;
  assign flit_address_o[7] = 1'b0;

  AND2X1 U6 ( .IN1(N19), .IN2(is_address), .Q(next_count[7]) );
  AND2X1 U7 ( .IN1(N18), .IN2(is_address), .Q(next_count[6]) );
  AND2X1 U9 ( .IN1(N17), .IN2(is_address), .Q(next_count[5]) );
  AND2X1 U10 ( .IN1(N16), .IN2(is_address), .Q(next_count[4]) );
  AND2X1 U11 ( .IN1(N15), .IN2(is_address), .Q(next_count[3]) );
  AND2X1 U12 ( .IN1(N14), .IN2(is_address), .Q(next_count[2]) );
  AND2X1 U13 ( .IN1(N13), .IN2(is_address), .Q(next_count[1]) );
  AND2X1 U14 ( .IN1(N12), .IN2(is_address), .Q(next_count[0]) );
  AND2X1 U16 ( .IN1(interface_flit_address[7]), .IN2(is_address), .Q(
        flit_address[7]) );
  AND2X1 U17 ( .IN1(interface_flit_address[6]), .IN2(is_address), .Q(
        flit_address[6]) );
  AND2X1 U18 ( .IN1(interface_flit_address[5]), .IN2(is_address), .Q(
        flit_address[5]) );
  AND2X1 U19 ( .IN1(interface_flit_address[4]), .IN2(is_address), .Q(
        flit_address[4]) );
  AND2X1 U20 ( .IN1(interface_flit_address[3]), .IN2(is_address), .Q(
        flit_address[3]) );
  AND2X1 U21 ( .IN1(interface_flit_address[2]), .IN2(is_address), .Q(
        flit_address[2]) );
  AND2X1 U22 ( .IN1(interface_flit_address[1]), .IN2(is_address), .Q(
        flit_address[1]) );
  AND2X1 U23 ( .IN1(interface_flit_address[0]), .IN2(is_address), .Q(
        flit_address[0]) );
  INVX0 U4 ( .INP(receiving_data), .ZN(n1) );
  NOR2X0 U5 ( .IN1(n1), .IN2(rst), .QN(is_address) );
  register_BITS8_0 count_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(next_count), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_8_0 address_reg ( .clk(clk), .enable_i(is_address), .reset(rst), 
        .data_i(flit_address), .data_o({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  address_counter_0_DW01_inc_0 r308 ( .A({1'b0, interface_flit_length}), .SUM(
        {SYNOPSYS_UNCONNECTED__0, N19, N18, N17, N16, N15, N14, N13, N12}) );
endmodule


module flipflop_BITS2_1 ( clk, data_i, data_o );
  input [1:0] data_i;
  output [1:0] data_o;
  input clk;


  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS2_1 ( clk, enable_i, reset, data_i, data_o );
  input [1:0] data_i;
  input [1:0] data_o;
  input clk, enable_i, reset;
  wire   n10, n11, n1, n5, n7, n8, n9;
  wire   [1:0] write_data;

  AOI22X1 U5 ( .IN1(enable_i), .IN2(data_i[1]), .IN3(n10), .IN4(n1), .QN(n9)
         );
  AOI22X1 U6 ( .IN1(data_i[0]), .IN2(enable_i), .IN3(n11), .IN4(n1), .QN(n8)
         );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n9), .QN(write_data[1]) );
  NOR2X0 U4 ( .IN1(reset), .IN2(n8), .QN(write_data[0]) );
  AND2X1 U7 ( .IN1(data_o[1]), .IN2(n7), .Q(n10) );
  AND2X1 U8 ( .IN1(data_o[0]), .IN2(n5), .Q(n11) );
  flipflop_BITS2_1 FF ( .clk(clk), .data_i(write_data), .data_o({n7, n5}) );
endmodule


module flipflop_BITS1_7 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_7 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_7 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter2_1 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [1:0] request;
  output [1:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   tail_en, n1, n2;
  wire   [1:0] req_i;
  wire   [1:0] req_o;

  AND3X1 U10 ( .IN1(request[1]), .IN2(n1), .IN3(n2), .Q(grant[1]) );
  AND3X1 U11 ( .IN1(request[0]), .IN2(n2), .IN3(request[1]), .Q(tail_en) );
  INVX0 U6 ( .INP(request[0]), .ZN(n1) );
  NOR2X0 U7 ( .IN1(buffer_full_i), .IN2(n1), .QN(grant[0]) );
  INVX0 U8 ( .INP(buffer_full_i), .ZN(n2) );
  OA21X1 U9 ( .IN1(request[1]), .IN2(request[0]), .IN3(n2), .Q(grant_v_o) );
  register_BITS2_1 req_record ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i({1'b1, 1'b0}), .data_o({1'b0, 1'b0}) );
  register_BITS1_7 tail ( .clk(clk), .enable_i(tail_en), .reset(rst), .data_i(
        1'b1), .data_o(1'b0) );
endmodule


module flipflop_BITS2_0 ( clk, data_i, data_o );
  input [1:0] data_i;
  output [1:0] data_o;
  input clk;


  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS2_0 ( clk, enable_i, reset, data_i, data_o );
  input [1:0] data_i;
  input [1:0] data_o;
  input clk, enable_i, reset;
  wire   n10, n11, n1, n5, n7, n8, n9;
  wire   [1:0] write_data;

  AOI22X1 U5 ( .IN1(enable_i), .IN2(data_i[1]), .IN3(n10), .IN4(n1), .QN(n9)
         );
  AOI22X1 U6 ( .IN1(data_i[0]), .IN2(enable_i), .IN3(n11), .IN4(n1), .QN(n8)
         );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n9), .QN(write_data[1]) );
  NOR2X0 U4 ( .IN1(reset), .IN2(n8), .QN(write_data[0]) );
  AND2X1 U7 ( .IN1(data_o[1]), .IN2(n7), .Q(n10) );
  AND2X1 U8 ( .IN1(data_o[0]), .IN2(n5), .Q(n11) );
  flipflop_BITS2_0 FF ( .clk(clk), .data_i(write_data), .data_o({n7, n5}) );
endmodule


module flipflop_BITS1_6 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_6 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_6 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter2_0 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [1:0] request;
  output [1:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   tail_en, n1, n2;
  wire   [1:0] req_i;
  wire   [1:0] req_o;

  AND3X1 U10 ( .IN1(request[1]), .IN2(n1), .IN3(n2), .Q(grant[1]) );
  AND3X1 U11 ( .IN1(request[0]), .IN2(n2), .IN3(request[1]), .Q(tail_en) );
  INVX0 U6 ( .INP(request[0]), .ZN(n1) );
  NOR2X0 U7 ( .IN1(buffer_full_i), .IN2(n1), .QN(grant[0]) );
  INVX0 U8 ( .INP(buffer_full_i), .ZN(n2) );
  OA21X1 U9 ( .IN1(request[1]), .IN2(request[0]), .IN3(n2), .Q(grant_v_o) );
  register_BITS2_0 req_record ( .clk(clk), .enable_i(tail_en), .reset(rst), 
        .data_i({1'b1, 1'b0}), .data_o({1'b0, 1'b0}) );
  register_BITS1_6 tail ( .clk(clk), .enable_i(tail_en), .reset(rst), .data_i(
        1'b1), .data_o(1'b0) );
endmodule


module flipflop_BITS4_8 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_8 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_8 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS4_7 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_7 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_7 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS4_6 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_6 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_6 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS1_5 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_5 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_5 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_4 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_4 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_4 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter4_2 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [3:0] request;
  output [3:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[2][3] , \req_i[2][2] , \req_i[2][1] , \req_i[2][0] ,
         \req_i[1][3] , \req_i[1][2] , \req_i[1][1] , \req_i[1][0] ,
         \req_i[0][3] , \req_i[0][2] , \req_i[0][1] , tail_en, N71, N265, N266,
         N267, N268, N276, N282, N291, N300, N301, N302, N303, n1, n2, n3, n4,
         n6, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21;
  wire   [2:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N265 = request[0];
  assign N266 = request[1];
  assign N267 = request[2];
  assign N268 = request[3];

  LATCHX1 shift_reg ( .CLK(1'b0), .D(1'b0), .Q(N71) );
  LATCHX1 \grant_reg[3]  ( .CLK(1'b1), .D(N303), .Q(grant[3]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N302), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N301), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N300), .Q(grant[0]) );
  LNANDX1 \req_i_reg[2][3]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][3] ) );
  LNANDX1 \req_i_reg[2][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][2] ) );
  LNANDX1 \req_i_reg[2][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][1] ) );
  LNANDX1 \req_i_reg[2][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][0] ) );
  LNANDX1 \req_i_reg[1][3]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][3] ) );
  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][3]  ( .CLK(tail_en), .D(N282), .Q(\req_i[0][3] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(n1), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(n4), .Q(\req_i[0][1] ) );
  LATCHX1 \tail_i_reg[0]  ( .CLK(tail_en), .D(N276), .Q(tail_i[0]) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N291), .D(tail_en), .Q(req_en[0]) );
  AND3X1 U35 ( .IN1(grant_v_o), .IN2(n19), .IN3(N267), .Q(N302) );
  NAND4X0 U37 ( .IN1(n17), .IN2(grant_v_o), .IN3(n16), .IN4(n20), .QN(N291) );
  AO21X1 U38 ( .IN1(n14), .IN2(n19), .IN3(buffer_full_i), .Q(n21) );
  NOR3X0 U39 ( .IN1(n4), .IN2(N282), .IN3(n1), .QN(n17) );
  NAND4X0 U41 ( .IN1(n11), .IN2(n13), .IN3(n9), .IN4(n10), .QN(N276) );
  AOI22X1 U42 ( .IN1(n2), .IN2(n15), .IN3(n15), .IN4(N265), .QN(n13) );
  AND2X1 U43 ( .IN1(N268), .IN2(n6), .Q(n15) );
  OA22X1 U44 ( .IN1(n6), .IN2(n18), .IN3(n6), .IN4(n3), .Q(n11) );
  INVX0 U15 ( .INP(N267), .ZN(n6) );
  INVX0 U16 ( .INP(n18), .ZN(n2) );
  NAND2X1 U17 ( .IN1(N266), .IN2(N265), .QN(n10) );
  NAND2X1 U18 ( .IN1(N267), .IN2(N268), .QN(n12) );
  INVX0 U19 ( .INP(N265), .ZN(n3) );
  NAND2X1 U20 ( .IN1(N266), .IN2(n3), .QN(n18) );
  NOR2X0 U21 ( .IN1(N266), .IN2(N265), .QN(n19) );
  INVX0 U22 ( .INP(n21), .ZN(grant_v_o) );
  NOR2X0 U23 ( .IN1(N268), .IN2(N267), .QN(n14) );
  NAND2X1 U24 ( .IN1(n15), .IN2(n19), .QN(n20) );
  NOR2X0 U25 ( .IN1(N265), .IN2(n2), .QN(n16) );
  NAND2X1 U26 ( .IN1(N71), .IN2(n7), .QN(n9) );
  INVX0 U27 ( .INP(n12), .ZN(n7) );
  INVX0 U28 ( .INP(n10), .ZN(n4) );
  INVX0 U29 ( .INP(n11), .ZN(n1) );
  NAND2X1 U30 ( .IN1(n13), .IN2(n12), .QN(N282) );
  NOR2X0 U31 ( .IN1(n21), .IN2(n17), .QN(tail_en) );
  NOR2X0 U32 ( .IN1(n3), .IN2(n21), .QN(N300) );
  NOR2X0 U33 ( .IN1(n18), .IN2(n21), .QN(N301) );
  NOR2X0 U34 ( .IN1(n21), .IN2(n20), .QN(N303) );
  register_BITS4_8 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][3] , \req_i[0][2] , \req_i[0][1] , 
        1'b0}), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS4_7 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][3] , \req_i[1][2] , \req_i[1][1] , 
        \req_i[1][0] }), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS4_6 \genblk1[2].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[2][3] , \req_i[2][2] , \req_i[2][1] , 
        \req_i[2][0] }), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS1_5 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(tail_i[0]), .data_o(1'b0) );
  register_BITS1_4 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module flipflop_BITS4_5 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_5 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_5 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS4_4 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_4 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_4 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS4_3 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_3 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_3 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS1_3 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_3 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_3 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_2 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_2 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_2 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter4_1 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [3:0] request;
  output [3:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[2][3] , \req_i[2][2] , \req_i[2][1] , \req_i[2][0] ,
         \req_i[1][3] , \req_i[1][2] , \req_i[1][1] , \req_i[1][0] ,
         \req_i[0][3] , \req_i[0][2] , \req_i[0][1] , tail_en, N71, N265, N266,
         N267, N268, N276, N282, N291, N300, N301, N302, N303, n1, n2, n3, n4,
         n6, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21;
  wire   [2:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N265 = request[0];
  assign N266 = request[1];
  assign N267 = request[2];
  assign N268 = request[3];

  LATCHX1 shift_reg ( .CLK(1'b0), .D(1'b0), .Q(N71) );
  LATCHX1 \grant_reg[3]  ( .CLK(1'b1), .D(N303), .Q(grant[3]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N302), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N301), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N300), .Q(grant[0]) );
  LNANDX1 \req_i_reg[2][3]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][3] ) );
  LNANDX1 \req_i_reg[2][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][2] ) );
  LNANDX1 \req_i_reg[2][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][1] ) );
  LNANDX1 \req_i_reg[2][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][0] ) );
  LNANDX1 \req_i_reg[1][3]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][3] ) );
  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][3]  ( .CLK(tail_en), .D(N282), .Q(\req_i[0][3] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(n1), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(n4), .Q(\req_i[0][1] ) );
  LATCHX1 \tail_i_reg[0]  ( .CLK(tail_en), .D(N276), .Q(tail_i[0]) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N291), .D(tail_en), .Q(req_en[0]) );
  AND3X1 U35 ( .IN1(grant_v_o), .IN2(n19), .IN3(N267), .Q(N302) );
  NAND4X0 U37 ( .IN1(n17), .IN2(grant_v_o), .IN3(n16), .IN4(n20), .QN(N291) );
  AO21X1 U38 ( .IN1(n14), .IN2(n19), .IN3(buffer_full_i), .Q(n21) );
  NOR3X0 U39 ( .IN1(n4), .IN2(N282), .IN3(n1), .QN(n17) );
  NAND4X0 U41 ( .IN1(n11), .IN2(n13), .IN3(n9), .IN4(n10), .QN(N276) );
  AOI22X1 U42 ( .IN1(n2), .IN2(n15), .IN3(n15), .IN4(N265), .QN(n13) );
  AND2X1 U43 ( .IN1(N268), .IN2(n6), .Q(n15) );
  OA22X1 U44 ( .IN1(n6), .IN2(n18), .IN3(n6), .IN4(n3), .Q(n11) );
  INVX0 U15 ( .INP(N267), .ZN(n6) );
  INVX0 U16 ( .INP(n18), .ZN(n2) );
  NAND2X1 U17 ( .IN1(N266), .IN2(N265), .QN(n10) );
  NAND2X1 U18 ( .IN1(N267), .IN2(N268), .QN(n12) );
  INVX0 U19 ( .INP(N265), .ZN(n3) );
  NAND2X1 U20 ( .IN1(N266), .IN2(n3), .QN(n18) );
  NOR2X0 U21 ( .IN1(N266), .IN2(N265), .QN(n19) );
  INVX0 U22 ( .INP(n21), .ZN(grant_v_o) );
  NOR2X0 U23 ( .IN1(N268), .IN2(N267), .QN(n14) );
  NAND2X1 U24 ( .IN1(n15), .IN2(n19), .QN(n20) );
  NOR2X0 U25 ( .IN1(N265), .IN2(n2), .QN(n16) );
  NAND2X1 U26 ( .IN1(N71), .IN2(n7), .QN(n9) );
  INVX0 U27 ( .INP(n12), .ZN(n7) );
  INVX0 U28 ( .INP(n10), .ZN(n4) );
  INVX0 U29 ( .INP(n11), .ZN(n1) );
  NAND2X1 U30 ( .IN1(n13), .IN2(n12), .QN(N282) );
  NOR2X0 U31 ( .IN1(n21), .IN2(n17), .QN(tail_en) );
  NOR2X0 U32 ( .IN1(n3), .IN2(n21), .QN(N300) );
  NOR2X0 U33 ( .IN1(n18), .IN2(n21), .QN(N301) );
  NOR2X0 U34 ( .IN1(n21), .IN2(n20), .QN(N303) );
  register_BITS4_5 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][3] , \req_i[0][2] , \req_i[0][1] , 
        1'b0}), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS4_4 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][3] , \req_i[1][2] , \req_i[1][1] , 
        \req_i[1][0] }), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS4_3 \genblk1[2].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[2][3] , \req_i[2][2] , \req_i[2][1] , 
        \req_i[2][0] }), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS1_3 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(tail_i[0]), .data_o(1'b0) );
  register_BITS1_2 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module flipflop_BITS4_2 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_2 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_2 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS4_1 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_1 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_1 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS4_0 ( clk, data_i, data_o );
  input [3:0] data_i;
  output [3:0] data_o;
  input clk;


  DFFX1 \data_o_reg[3]  ( .D(data_i[3]), .CLK(clk), .Q(data_o[3]) );
  DFFX1 \data_o_reg[2]  ( .D(data_i[2]), .CLK(clk), .Q(data_o[2]) );
  DFFX1 \data_o_reg[1]  ( .D(data_i[1]), .CLK(clk), .Q(data_o[1]) );
  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS4_0 ( clk, enable_i, reset, data_i, data_o );
  input [3:0] data_i;
  input [3:0] data_o;
  input clk, enable_i, reset;
  wire   n14, n15, n16, n17, n1, n5, n7, n9, n11, n12, n13;
  wire   [3:0] write_data;

  AO22X1 U5 ( .IN1(data_i[3]), .IN2(n13), .IN3(n14), .IN4(n12), .Q(
        write_data[3]) );
  AO22X1 U6 ( .IN1(data_i[2]), .IN2(n13), .IN3(n15), .IN4(n12), .Q(
        write_data[2]) );
  AO22X1 U7 ( .IN1(data_i[1]), .IN2(n13), .IN3(n16), .IN4(n12), .Q(
        write_data[1]) );
  AO22X1 U8 ( .IN1(data_i[0]), .IN2(n13), .IN3(n17), .IN4(n12), .Q(
        write_data[0]) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(enable_i), .IN2(reset), .QN(n12) );
  NOR2X0 U4 ( .IN1(n1), .IN2(reset), .QN(n13) );
  AND2X1 U9 ( .IN1(data_o[3]), .IN2(n11), .Q(n14) );
  AND2X1 U10 ( .IN1(data_o[2]), .IN2(n9), .Q(n15) );
  AND2X1 U11 ( .IN1(data_o[1]), .IN2(n7), .Q(n16) );
  AND2X1 U12 ( .IN1(data_o[0]), .IN2(n5), .Q(n17) );
  flipflop_BITS4_0 FF ( .clk(clk), .data_i(write_data), .data_o({n11, n9, n7, 
        n5}) );
endmodule


module flipflop_BITS1_1 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_1 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_1 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module flipflop_BITS1_0 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  DFFX1 \data_o_reg[0]  ( .D(data_i[0]), .CLK(clk), .Q(data_o[0]) );
endmodule


module register_BITS1_0 ( clk, enable_i, reset, data_i, data_o );
  input [0:0] data_i;
  input [0:0] data_o;
  input clk, enable_i, reset;
  wire   n6, \write_data[0] , n1, n4, n5;

  AOI22X1 U4 ( .IN1(enable_i), .IN2(data_i[0]), .IN3(n6), .IN4(n1), .QN(n5) );
  INVX0 U2 ( .INP(enable_i), .ZN(n1) );
  NOR2X0 U3 ( .IN1(reset), .IN2(n5), .QN(\write_data[0] ) );
  AND2X1 U5 ( .IN1(data_o[0]), .IN2(n4), .Q(n6) );
  flipflop_BITS1_0 FF ( .clk(clk), .data_i(\write_data[0] ), .data_o(n4) );
endmodule


module arbiter4_0 ( clk, rst, request, buffer_full_i, grant, grant_v_o );
  input [3:0] request;
  output [3:0] grant;
  input clk, rst, buffer_full_i;
  output grant_v_o;
  wire   \req_i[2][3] , \req_i[2][2] , \req_i[2][1] , \req_i[2][0] ,
         \req_i[1][3] , \req_i[1][2] , \req_i[1][1] , \req_i[1][0] ,
         \req_i[0][3] , \req_i[0][2] , \req_i[0][1] , tail_en, N71, N265, N266,
         N267, N268, N276, N282, N291, N300, N301, N302, N303, n1, n2, n3, n4,
         n6, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21;
  wire   [2:0] req_en;
  wire   [1:0] tail_i;
  wire   [1:0] tail_o;
  assign N265 = request[0];
  assign N266 = request[1];
  assign N267 = request[2];
  assign N268 = request[3];

  LATCHX1 shift_reg ( .CLK(1'b0), .D(1'b0), .Q(N71) );
  LATCHX1 \grant_reg[3]  ( .CLK(1'b1), .D(N303), .Q(grant[3]) );
  LATCHX1 \grant_reg[2]  ( .CLK(1'b1), .D(N302), .Q(grant[2]) );
  LATCHX1 \grant_reg[1]  ( .CLK(1'b1), .D(N301), .Q(grant[1]) );
  LATCHX1 \grant_reg[0]  ( .CLK(1'b1), .D(N300), .Q(grant[0]) );
  LNANDX1 \req_i_reg[2][3]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][3] ) );
  LNANDX1 \req_i_reg[2][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][2] ) );
  LNANDX1 \req_i_reg[2][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][1] ) );
  LNANDX1 \req_i_reg[2][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[2][0] ) );
  LNANDX1 \req_i_reg[1][3]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][3] ) );
  LNANDX1 \req_i_reg[1][2]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][2] ) );
  LNANDX1 \req_i_reg[1][1]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][1] ) );
  LNANDX1 \req_i_reg[1][0]  ( .RIN(1'b1), .SIN(1'b1), .Q(\req_i[1][0] ) );
  LATCHX1 \req_i_reg[0][3]  ( .CLK(tail_en), .D(N282), .Q(\req_i[0][3] ) );
  LATCHX1 \req_i_reg[0][2]  ( .CLK(tail_en), .D(n1), .Q(\req_i[0][2] ) );
  LATCHX1 \req_i_reg[0][1]  ( .CLK(tail_en), .D(n4), .Q(\req_i[0][1] ) );
  LATCHX1 \tail_i_reg[0]  ( .CLK(tail_en), .D(N276), .Q(tail_i[0]) );
  LATCHX1 \req_en_reg[0]  ( .CLK(N291), .D(tail_en), .Q(req_en[0]) );
  AND3X1 U35 ( .IN1(grant_v_o), .IN2(n19), .IN3(N267), .Q(N302) );
  NAND4X0 U37 ( .IN1(n17), .IN2(grant_v_o), .IN3(n16), .IN4(n20), .QN(N291) );
  AO21X1 U38 ( .IN1(n14), .IN2(n19), .IN3(buffer_full_i), .Q(n21) );
  NOR3X0 U39 ( .IN1(n4), .IN2(N282), .IN3(n1), .QN(n17) );
  NAND4X0 U41 ( .IN1(n11), .IN2(n13), .IN3(n9), .IN4(n10), .QN(N276) );
  AOI22X1 U42 ( .IN1(n2), .IN2(n15), .IN3(n15), .IN4(N265), .QN(n13) );
  AND2X1 U43 ( .IN1(N268), .IN2(n6), .Q(n15) );
  OA22X1 U44 ( .IN1(n6), .IN2(n18), .IN3(n6), .IN4(n3), .Q(n11) );
  INVX0 U15 ( .INP(N267), .ZN(n6) );
  INVX0 U16 ( .INP(n18), .ZN(n2) );
  NAND2X1 U17 ( .IN1(N266), .IN2(N265), .QN(n10) );
  NAND2X1 U18 ( .IN1(N267), .IN2(N268), .QN(n12) );
  INVX0 U19 ( .INP(N265), .ZN(n3) );
  NAND2X1 U20 ( .IN1(N266), .IN2(n3), .QN(n18) );
  NOR2X0 U21 ( .IN1(N266), .IN2(N265), .QN(n19) );
  INVX0 U22 ( .INP(n21), .ZN(grant_v_o) );
  NOR2X0 U23 ( .IN1(N268), .IN2(N267), .QN(n14) );
  NAND2X1 U24 ( .IN1(n15), .IN2(n19), .QN(n20) );
  NOR2X0 U25 ( .IN1(N265), .IN2(n2), .QN(n16) );
  NAND2X1 U26 ( .IN1(N71), .IN2(n7), .QN(n9) );
  INVX0 U27 ( .INP(n12), .ZN(n7) );
  INVX0 U28 ( .INP(n10), .ZN(n4) );
  INVX0 U29 ( .INP(n11), .ZN(n1) );
  NAND2X1 U30 ( .IN1(n13), .IN2(n12), .QN(N282) );
  NOR2X0 U31 ( .IN1(n21), .IN2(n17), .QN(tail_en) );
  NOR2X0 U32 ( .IN1(n3), .IN2(n21), .QN(N300) );
  NOR2X0 U33 ( .IN1(n18), .IN2(n21), .QN(N301) );
  NOR2X0 U34 ( .IN1(n21), .IN2(n20), .QN(N303) );
  register_BITS4_2 \genblk1[0].req_record  ( .clk(clk), .enable_i(req_en[0]), 
        .reset(rst), .data_i({\req_i[0][3] , \req_i[0][2] , \req_i[0][1] , 
        1'b0}), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS4_1 \genblk1[1].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[1][3] , \req_i[1][2] , \req_i[1][1] , 
        \req_i[1][0] }), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS4_0 \genblk1[2].req_record  ( .clk(clk), .enable_i(1'b0), 
        .reset(rst), .data_i({\req_i[2][3] , \req_i[2][2] , \req_i[2][1] , 
        \req_i[2][0] }), .data_o({1'b0, 1'b0, 1'b0, 1'b0}) );
  register_BITS1_1 \genblk2[0].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(tail_i[0]), .data_o(1'b0) );
  register_BITS1_0 \genblk2[1].tail  ( .clk(clk), .enable_i(tail_en), .reset(
        rst), .data_i(1'b0), .data_o(1'b0) );
endmodule


module dccl_4 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_3 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_2 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_1 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module dccl_0 ( packet_addr_y_i, packet_addr_x_i, local_addr_y_i, 
        local_addr_x_i, packet_valid_i, north_req, east_req, south_req, 
        west_req, local_req );
  input [3:0] packet_addr_y_i;
  input [3:0] packet_addr_x_i;
  input [3:0] local_addr_y_i;
  input [3:0] local_addr_x_i;
  input packet_valid_i;
  output north_req, east_req, south_req, west_req, local_req;
  wire   N18, N20, N21, N22, N23, n1, n2, n3, n4, n5, n6, n7, n8, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  LATCHX1 north_req_reg ( .CLK(1'b1), .D(N20), .Q(north_req) );
  LATCHX1 east_req_reg ( .CLK(1'b1), .D(N21), .Q(east_req) );
  LATCHX1 south_req_reg ( .CLK(1'b1), .D(N22), .Q(south_req) );
  LATCHX1 west_req_reg ( .CLK(1'b1), .D(N23), .Q(west_req) );
  LATCHX1 local_req_reg ( .CLK(1'b1), .D(N18), .Q(local_req) );
  AND3X1 U26 ( .IN1(n1), .IN2(n62), .IN3(n2), .Q(N23) );
  NOR3X0 U27 ( .IN1(n62), .IN2(n59), .IN3(n61), .QN(N21) );
  AO22X1 U28 ( .IN1(local_addr_x_i[3]), .IN2(n58), .IN3(n57), .IN4(n14), .Q(
        n62) );
  OR2X1 U29 ( .IN1(n58), .IN2(local_addr_x_i[3]), .Q(n57) );
  AO22X1 U30 ( .IN1(local_addr_x_i[2]), .IN2(n8), .IN3(n56), .IN4(n55), .Q(n58) );
  AO21X1 U31 ( .IN1(local_addr_x_i[1]), .IN2(n7), .IN3(local_addr_x_i[0]), .Q(
        n55) );
  AND3X1 U32 ( .IN1(n1), .IN2(n59), .IN3(n60), .Q(N20) );
  AO22X1 U33 ( .IN1(local_addr_y_i[3]), .IN2(n52), .IN3(n51), .IN4(n6), .Q(n60) );
  OR2X1 U34 ( .IN1(n52), .IN2(local_addr_y_i[3]), .Q(n51) );
  AO22X1 U35 ( .IN1(local_addr_y_i[2]), .IN2(n4), .IN3(n50), .IN4(n49), .Q(n52) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n16), .IN3(packet_addr_y_i[0]), .QN(n49) );
  NAND4X0 U38 ( .IN1(n25), .IN2(n2), .IN3(n24), .IN4(n23), .QN(n45) );
  AOI221X1 U39 ( .IN1(n8), .IN2(local_addr_x_i[2]), .IN3(n7), .IN4(
        local_addr_x_i[1]), .IN5(n22), .QN(n23) );
  OR2X1 U40 ( .IN1(n54), .IN2(n53), .Q(n22) );
  XNOR2X1 U41 ( .IN1(local_addr_x_i[0]), .IN2(packet_addr_x_i[0]), .Q(n24) );
  NAND4X0 U42 ( .IN1(n21), .IN2(n20), .IN3(n19), .IN4(n46), .QN(n59) );
  AOI21X1 U43 ( .IN1(n3), .IN2(local_addr_y_i[1]), .IN3(n47), .QN(n19) );
  XOR2X1 U44 ( .IN1(n16), .IN2(packet_addr_y_i[0]), .Q(n20) );
  XOR2X1 U45 ( .IN1(local_addr_y_i[3]), .IN2(n6), .Q(n18) );
  XOR2X1 U46 ( .IN1(local_addr_x_i[3]), .IN2(n14), .Q(n25) );
  NOR2X0 U3 ( .IN1(n7), .IN2(local_addr_x_i[1]), .QN(n53) );
  NOR2X0 U4 ( .IN1(n8), .IN2(local_addr_x_i[2]), .QN(n54) );
  INVX0 U5 ( .INP(packet_addr_x_i[3]), .ZN(n14) );
  INVX0 U6 ( .INP(packet_addr_x_i[1]), .ZN(n7) );
  NOR2X0 U7 ( .IN1(n54), .IN2(n53), .QN(n56) );
  INVX0 U8 ( .INP(packet_addr_x_i[2]), .ZN(n8) );
  INVX0 U9 ( .INP(packet_addr_y_i[1]), .ZN(n3) );
  NOR2X0 U10 ( .IN1(n3), .IN2(local_addr_y_i[1]), .QN(n47) );
  INVX0 U11 ( .INP(local_addr_y_i[2]), .ZN(n17) );
  INVX0 U12 ( .INP(local_addr_y_i[0]), .ZN(n16) );
  NAND2X1 U13 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .QN(n46) );
  INVX0 U14 ( .INP(packet_addr_y_i[3]), .ZN(n6) );
  NAND2X1 U15 ( .IN1(local_addr_y_i[1]), .IN2(n3), .QN(n48) );
  NOR2X0 U16 ( .IN1(n47), .IN2(n5), .QN(n50) );
  INVX0 U17 ( .INP(n46), .ZN(n5) );
  INVX0 U18 ( .INP(n59), .ZN(n2) );
  NAND2X1 U19 ( .IN1(packet_valid_i), .IN2(n45), .QN(n61) );
  OA21X1 U20 ( .IN1(packet_addr_y_i[2]), .IN2(n17), .IN3(n18), .Q(n21) );
  INVX0 U21 ( .INP(packet_addr_y_i[2]), .ZN(n4) );
  INVX0 U22 ( .INP(n61), .ZN(n1) );
  NOR2X0 U23 ( .IN1(n15), .IN2(n45), .QN(N18) );
  INVX0 U24 ( .INP(packet_valid_i), .ZN(n15) );
  NOR2X0 U25 ( .IN1(n61), .IN2(n60), .QN(N22) );
endmodule


module controller5_0 ( clk, rst, .packet_addr({\packet_addr[4][7] , 
        \packet_addr[4][6] , \packet_addr[4][5] , \packet_addr[4][4] , 
        \packet_addr[4][3] , \packet_addr[4][2] , \packet_addr[4][1] , 
        \packet_addr[4][0] , \packet_addr[3][7] , \packet_addr[3][6] , 
        \packet_addr[3][5] , \packet_addr[3][4] , \packet_addr[3][3] , 
        \packet_addr[3][2] , \packet_addr[3][1] , \packet_addr[3][0] , 
        \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] , 
        \packet_addr[2][4] , \packet_addr[2][3] , \packet_addr[2][2] , 
        \packet_addr[2][1] , \packet_addr[2][0] , \packet_addr[1][7] , 
        \packet_addr[1][6] , \packet_addr[1][5] , \packet_addr[1][4] , 
        \packet_addr[1][3] , \packet_addr[1][2] , \packet_addr[1][1] , 
        \packet_addr[1][0] , \packet_addr[0][7] , \packet_addr[0][6] , 
        \packet_addr[0][5] , \packet_addr[0][4] , \packet_addr[0][3] , 
        \packet_addr[0][2] , \packet_addr[0][1] , \packet_addr[0][0] }), 
        local_addr, packet_valid, buffer_full_in, grant_0, grant_1, grant_2, 
        grant_3, grant_4, grant_v, pop_v );
  input [7:0] local_addr;
  input [4:0] packet_valid;
  input [4:0] buffer_full_in;
  output [1:0] grant_0;
  output [1:0] grant_1;
  output [3:0] grant_2;
  output [3:0] grant_3;
  output [3:0] grant_4;
  output [4:0] grant_v;
  output [4:0] pop_v;
  input clk, rst, \packet_addr[4][7] , \packet_addr[4][6] ,
         \packet_addr[4][5] , \packet_addr[4][4] , \packet_addr[4][3] ,
         \packet_addr[4][2] , \packet_addr[4][1] , \packet_addr[4][0] ,
         \packet_addr[3][7] , \packet_addr[3][6] , \packet_addr[3][5] ,
         \packet_addr[3][4] , \packet_addr[3][3] , \packet_addr[3][2] ,
         \packet_addr[3][1] , \packet_addr[3][0] , \packet_addr[2][7] ,
         \packet_addr[2][6] , \packet_addr[2][5] , \packet_addr[2][4] ,
         \packet_addr[2][3] , \packet_addr[2][2] , \packet_addr[2][1] ,
         \packet_addr[2][0] , \packet_addr[1][7] , \packet_addr[1][6] ,
         \packet_addr[1][5] , \packet_addr[1][4] , \packet_addr[1][3] ,
         \packet_addr[1][2] , \packet_addr[1][1] , \packet_addr[1][0] ,
         \packet_addr[0][7] , \packet_addr[0][6] , \packet_addr[0][5] ,
         \packet_addr[0][4] , \packet_addr[0][3] , \packet_addr[0][2] ,
         \packet_addr[0][1] , \packet_addr[0][0] ;
  wire   \request[4][3] , \request[4][2] , \request[4][1] , \request[4][0] ,
         \request[3][3] , \request[3][2] , \request[3][1] , \request[3][0] ,
         \request[2][3] , \request[2][2] , \request[2][1] , \request[2][0] ,
         \request[1][1] , \request[1][0] , \request[0][1] , \request[0][0] ;

  OR4X1 U1 ( .IN1(grant_1[1]), .IN2(grant_0[1]), .IN3(grant_3[3]), .IN4(
        grant_2[3]), .Q(pop_v[4]) );
  OR2X1 U2 ( .IN1(grant_2[2]), .IN2(grant_4[3]), .Q(pop_v[3]) );
  OR2X1 U3 ( .IN1(grant_3[2]), .IN2(grant_4[2]), .Q(pop_v[2]) );
  OR4X1 U4 ( .IN1(grant_2[1]), .IN2(grant_0[0]), .IN3(grant_4[1]), .IN4(
        grant_3[1]), .Q(pop_v[1]) );
  OR4X1 U5 ( .IN1(grant_2[0]), .IN2(grant_1[0]), .IN3(grant_4[0]), .IN4(
        grant_3[0]), .Q(pop_v[0]) );
  arbiter2_1 arbiter_n ( .clk(clk), .rst(rst), .request({\request[0][1] , 
        \request[0][0] }), .buffer_full_i(buffer_full_in[0]), .grant(grant_0), 
        .grant_v_o(grant_v[0]) );
  arbiter2_0 arbiter_s ( .clk(clk), .rst(rst), .request({\request[1][1] , 
        \request[1][0] }), .buffer_full_i(buffer_full_in[1]), .grant(grant_1), 
        .grant_v_o(grant_v[1]) );
  arbiter4_2 arbiter_e ( .clk(clk), .rst(rst), .request({\request[2][3] , 
        \request[2][2] , \request[2][1] , \request[2][0] }), .buffer_full_i(
        buffer_full_in[2]), .grant(grant_2), .grant_v_o(grant_v[2]) );
  arbiter4_1 arbiter_w ( .clk(clk), .rst(rst), .request({\request[3][3] , 
        \request[3][2] , \request[3][1] , \request[3][0] }), .buffer_full_i(
        buffer_full_in[3]), .grant(grant_3), .grant_v_o(grant_v[3]) );
  arbiter4_0 arbiter_l ( .clk(clk), .rst(rst), .request({\request[4][3] , 
        \request[4][2] , \request[4][1] , \request[4][0] }), .buffer_full_i(
        buffer_full_in[4]), .grant(grant_4), .grant_v_o(grant_v[4]) );
  dccl_4 dccl_n ( .packet_addr_y_i({\packet_addr[0][3] , \packet_addr[0][2] , 
        \packet_addr[0][1] , \packet_addr[0][0] }), .packet_addr_x_i({
        \packet_addr[0][7] , \packet_addr[0][6] , \packet_addr[0][5] , 
        \packet_addr[0][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[0]), 
        .east_req(\request[2][0] ), .south_req(\request[1][0] ), .west_req(
        \request[3][0] ), .local_req(\request[4][0] ) );
  dccl_3 dccl_s ( .packet_addr_y_i({\packet_addr[1][3] , \packet_addr[1][2] , 
        \packet_addr[1][1] , \packet_addr[1][0] }), .packet_addr_x_i({
        \packet_addr[1][7] , \packet_addr[1][6] , \packet_addr[1][5] , 
        \packet_addr[1][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[1]), 
        .north_req(\request[0][0] ), .east_req(\request[2][1] ), .west_req(
        \request[3][1] ), .local_req(\request[4][1] ) );
  dccl_2 dccl_e ( .packet_addr_y_i({\packet_addr[2][3] , \packet_addr[2][2] , 
        \packet_addr[2][1] , \packet_addr[2][0] }), .packet_addr_x_i({
        \packet_addr[2][7] , \packet_addr[2][6] , \packet_addr[2][5] , 
        \packet_addr[2][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[2]), 
        .west_req(\request[3][2] ), .local_req(\request[4][2] ) );
  dccl_1 dccl_w ( .packet_addr_y_i({\packet_addr[3][3] , \packet_addr[3][2] , 
        \packet_addr[3][1] , \packet_addr[3][0] }), .packet_addr_x_i({
        \packet_addr[3][7] , \packet_addr[3][6] , \packet_addr[3][5] , 
        \packet_addr[3][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[3]), 
        .east_req(\request[2][2] ), .local_req(\request[4][3] ) );
  dccl_0 dccl_l ( .packet_addr_y_i({\packet_addr[4][3] , \packet_addr[4][2] , 
        \packet_addr[4][1] , \packet_addr[4][0] }), .packet_addr_x_i({
        \packet_addr[4][7] , \packet_addr[4][6] , \packet_addr[4][5] , 
        \packet_addr[4][4] }), .local_addr_y_i(local_addr[3:0]), 
        .local_addr_x_i(local_addr[7:4]), .packet_valid_i(packet_valid[4]), 
        .north_req(\request[0][1] ), .east_req(\request[2][3] ), .south_req(
        \request[1][1] ), .west_req(\request[3][3] ) );
endmodule


module mux2_1_1 ( data0, data1, select0, select1, data_o );
  input [15:0] data0;
  input [15:0] data1;
  output [15:0] data_o;
  input select0, select1;
  wire   n1, n4, n5;

  AO22X1 U4 ( .IN1(data1[9]), .IN2(n5), .IN3(data0[9]), .IN4(n4), .Q(data_o[9]) );
  AO22X1 U5 ( .IN1(data1[8]), .IN2(n5), .IN3(data0[8]), .IN4(n4), .Q(data_o[8]) );
  AO22X1 U6 ( .IN1(data1[7]), .IN2(n5), .IN3(data0[7]), .IN4(n4), .Q(data_o[7]) );
  AO22X1 U7 ( .IN1(data1[6]), .IN2(n5), .IN3(data0[6]), .IN4(n4), .Q(data_o[6]) );
  AO22X1 U8 ( .IN1(data1[5]), .IN2(n5), .IN3(data0[5]), .IN4(n4), .Q(data_o[5]) );
  AO22X1 U9 ( .IN1(data1[4]), .IN2(n5), .IN3(data0[4]), .IN4(n4), .Q(data_o[4]) );
  AO22X1 U10 ( .IN1(data1[3]), .IN2(n5), .IN3(data0[3]), .IN4(n4), .Q(
        data_o[3]) );
  AO22X1 U11 ( .IN1(data1[2]), .IN2(n5), .IN3(data0[2]), .IN4(n4), .Q(
        data_o[2]) );
  AO22X1 U12 ( .IN1(data1[1]), .IN2(n5), .IN3(data0[1]), .IN4(n4), .Q(
        data_o[1]) );
  AO22X1 U13 ( .IN1(data1[15]), .IN2(n5), .IN3(data0[15]), .IN4(n4), .Q(
        data_o[15]) );
  AO22X1 U14 ( .IN1(data1[14]), .IN2(n5), .IN3(data0[14]), .IN4(n4), .Q(
        data_o[14]) );
  AO22X1 U15 ( .IN1(data1[13]), .IN2(n5), .IN3(data0[13]), .IN4(n4), .Q(
        data_o[13]) );
  AO22X1 U16 ( .IN1(data1[12]), .IN2(n5), .IN3(data0[12]), .IN4(n4), .Q(
        data_o[12]) );
  AO22X1 U17 ( .IN1(data1[11]), .IN2(n5), .IN3(data0[11]), .IN4(n4), .Q(
        data_o[11]) );
  AO22X1 U18 ( .IN1(data1[10]), .IN2(n5), .IN3(data0[10]), .IN4(n4), .Q(
        data_o[10]) );
  AO22X1 U19 ( .IN1(data1[0]), .IN2(n5), .IN3(data0[0]), .IN4(n4), .Q(
        data_o[0]) );
  INVX0 U2 ( .INP(select1), .ZN(n1) );
  AND2X1 U3 ( .IN1(select0), .IN2(n1), .Q(n4) );
  NOR2X0 U20 ( .IN1(n1), .IN2(select0), .QN(n5) );
endmodule


module mux2_1_0 ( data0, data1, select0, select1, data_o );
  input [15:0] data0;
  input [15:0] data1;
  output [15:0] data_o;
  input select0, select1;
  wire   n1, n4, n5;

  AO22X1 U4 ( .IN1(data1[9]), .IN2(n5), .IN3(data0[9]), .IN4(n4), .Q(data_o[9]) );
  AO22X1 U5 ( .IN1(data1[8]), .IN2(n5), .IN3(data0[8]), .IN4(n4), .Q(data_o[8]) );
  AO22X1 U6 ( .IN1(data1[7]), .IN2(n5), .IN3(data0[7]), .IN4(n4), .Q(data_o[7]) );
  AO22X1 U7 ( .IN1(data1[6]), .IN2(n5), .IN3(data0[6]), .IN4(n4), .Q(data_o[6]) );
  AO22X1 U8 ( .IN1(data1[5]), .IN2(n5), .IN3(data0[5]), .IN4(n4), .Q(data_o[5]) );
  AO22X1 U9 ( .IN1(data1[4]), .IN2(n5), .IN3(data0[4]), .IN4(n4), .Q(data_o[4]) );
  AO22X1 U10 ( .IN1(data1[3]), .IN2(n5), .IN3(data0[3]), .IN4(n4), .Q(
        data_o[3]) );
  AO22X1 U11 ( .IN1(data1[2]), .IN2(n5), .IN3(data0[2]), .IN4(n4), .Q(
        data_o[2]) );
  AO22X1 U12 ( .IN1(data1[1]), .IN2(n5), .IN3(data0[1]), .IN4(n4), .Q(
        data_o[1]) );
  AO22X1 U13 ( .IN1(data1[15]), .IN2(n5), .IN3(data0[15]), .IN4(n4), .Q(
        data_o[15]) );
  AO22X1 U14 ( .IN1(data1[14]), .IN2(n5), .IN3(data0[14]), .IN4(n4), .Q(
        data_o[14]) );
  AO22X1 U15 ( .IN1(data1[13]), .IN2(n5), .IN3(data0[13]), .IN4(n4), .Q(
        data_o[13]) );
  AO22X1 U16 ( .IN1(data1[12]), .IN2(n5), .IN3(data0[12]), .IN4(n4), .Q(
        data_o[12]) );
  AO22X1 U17 ( .IN1(data1[11]), .IN2(n5), .IN3(data0[11]), .IN4(n4), .Q(
        data_o[11]) );
  AO22X1 U18 ( .IN1(data1[10]), .IN2(n5), .IN3(data0[10]), .IN4(n4), .Q(
        data_o[10]) );
  AO22X1 U19 ( .IN1(data1[0]), .IN2(n5), .IN3(data0[0]), .IN4(n4), .Q(
        data_o[0]) );
  INVX0 U2 ( .INP(select1), .ZN(n1) );
  AND2X1 U3 ( .IN1(select0), .IN2(n1), .Q(n4) );
  NOR2X0 U20 ( .IN1(n1), .IN2(select0), .QN(n5) );
endmodule


module mux4_1_2 ( data0, data1, data2, data3, select0, select1, select2, 
        select3, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  input [15:0] data3;
  output [15:0] data_o;
  input select0, select1, select2, select3;
  wire   n1, n2, n3, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43;

  AO221X1 U5 ( .IN1(data1[9]), .IN2(n43), .IN3(data0[9]), .IN4(n42), .IN5(n41), 
        .Q(data_o[9]) );
  AO22X1 U6 ( .IN1(data2[9]), .IN2(n40), .IN3(data3[9]), .IN4(n39), .Q(n41) );
  AO221X1 U7 ( .IN1(data1[8]), .IN2(n43), .IN3(data0[8]), .IN4(n42), .IN5(n38), 
        .Q(data_o[8]) );
  AO22X1 U8 ( .IN1(data2[8]), .IN2(n40), .IN3(data3[8]), .IN4(n39), .Q(n38) );
  AO221X1 U9 ( .IN1(data1[7]), .IN2(n43), .IN3(data0[7]), .IN4(n42), .IN5(n37), 
        .Q(data_o[7]) );
  AO22X1 U10 ( .IN1(data2[7]), .IN2(n40), .IN3(data3[7]), .IN4(n39), .Q(n37)
         );
  AO221X1 U11 ( .IN1(data1[6]), .IN2(n43), .IN3(data0[6]), .IN4(n42), .IN5(n36), .Q(data_o[6]) );
  AO22X1 U12 ( .IN1(data2[6]), .IN2(n40), .IN3(data3[6]), .IN4(n39), .Q(n36)
         );
  AO221X1 U13 ( .IN1(data1[5]), .IN2(n43), .IN3(data0[5]), .IN4(n42), .IN5(n35), .Q(data_o[5]) );
  AO22X1 U14 ( .IN1(data2[5]), .IN2(n40), .IN3(data3[5]), .IN4(n39), .Q(n35)
         );
  AO221X1 U15 ( .IN1(data1[4]), .IN2(n43), .IN3(data0[4]), .IN4(n42), .IN5(n34), .Q(data_o[4]) );
  AO22X1 U16 ( .IN1(data2[4]), .IN2(n40), .IN3(data3[4]), .IN4(n39), .Q(n34)
         );
  AO221X1 U17 ( .IN1(data1[3]), .IN2(n43), .IN3(data0[3]), .IN4(n42), .IN5(n33), .Q(data_o[3]) );
  AO22X1 U18 ( .IN1(data2[3]), .IN2(n40), .IN3(data3[3]), .IN4(n39), .Q(n33)
         );
  AO221X1 U19 ( .IN1(data1[2]), .IN2(n43), .IN3(data0[2]), .IN4(n42), .IN5(n32), .Q(data_o[2]) );
  AO22X1 U20 ( .IN1(data2[2]), .IN2(n40), .IN3(data3[2]), .IN4(n39), .Q(n32)
         );
  AO221X1 U21 ( .IN1(data1[1]), .IN2(n43), .IN3(data0[1]), .IN4(n42), .IN5(n31), .Q(data_o[1]) );
  AO22X1 U22 ( .IN1(data2[1]), .IN2(n40), .IN3(data3[1]), .IN4(n39), .Q(n31)
         );
  AO221X1 U23 ( .IN1(data1[15]), .IN2(n43), .IN3(data0[15]), .IN4(n42), .IN5(
        n30), .Q(data_o[15]) );
  AO22X1 U24 ( .IN1(data2[15]), .IN2(n40), .IN3(data3[15]), .IN4(n39), .Q(n30)
         );
  AO221X1 U25 ( .IN1(data1[14]), .IN2(n43), .IN3(data0[14]), .IN4(n42), .IN5(
        n29), .Q(data_o[14]) );
  AO22X1 U26 ( .IN1(data2[14]), .IN2(n40), .IN3(data3[14]), .IN4(n39), .Q(n29)
         );
  AO221X1 U27 ( .IN1(data1[13]), .IN2(n43), .IN3(data0[13]), .IN4(n42), .IN5(
        n28), .Q(data_o[13]) );
  AO22X1 U28 ( .IN1(data2[13]), .IN2(n40), .IN3(data3[13]), .IN4(n39), .Q(n28)
         );
  AO221X1 U29 ( .IN1(data1[12]), .IN2(n43), .IN3(data0[12]), .IN4(n42), .IN5(
        n27), .Q(data_o[12]) );
  AO22X1 U30 ( .IN1(data2[12]), .IN2(n40), .IN3(data3[12]), .IN4(n39), .Q(n27)
         );
  AO221X1 U31 ( .IN1(data1[11]), .IN2(n43), .IN3(data0[11]), .IN4(n42), .IN5(
        n26), .Q(data_o[11]) );
  AO22X1 U32 ( .IN1(data2[11]), .IN2(n40), .IN3(data3[11]), .IN4(n39), .Q(n26)
         );
  AO221X1 U33 ( .IN1(data1[10]), .IN2(n43), .IN3(data0[10]), .IN4(n42), .IN5(
        n25), .Q(data_o[10]) );
  AO22X1 U34 ( .IN1(data2[10]), .IN2(n40), .IN3(data3[10]), .IN4(n39), .Q(n25)
         );
  AO221X1 U35 ( .IN1(data1[0]), .IN2(n43), .IN3(data0[0]), .IN4(n42), .IN5(n24), .Q(data_o[0]) );
  AO22X1 U36 ( .IN1(data2[0]), .IN2(n40), .IN3(data3[0]), .IN4(n39), .Q(n24)
         );
  INVX0 U2 ( .INP(select2), .ZN(n1) );
  NOR4X0 U3 ( .IN1(n1), .IN2(select0), .IN3(select1), .IN4(select3), .QN(n40)
         );
  AND4X1 U4 ( .IN1(select3), .IN2(n3), .IN3(n2), .IN4(n1), .Q(n39) );
  INVX0 U37 ( .INP(select0), .ZN(n3) );
  INVX0 U38 ( .INP(select1), .ZN(n2) );
  NOR4X0 U39 ( .IN1(n3), .IN2(select1), .IN3(select2), .IN4(select3), .QN(n42)
         );
  NOR4X0 U40 ( .IN1(n2), .IN2(select0), .IN3(select2), .IN4(select3), .QN(n43)
         );
endmodule


module mux4_1_1 ( data0, data1, data2, data3, select0, select1, select2, 
        select3, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  input [15:0] data3;
  output [15:0] data_o;
  input select0, select1, select2, select3;
  wire   n1, n2, n3, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43;

  AO221X1 U5 ( .IN1(data1[9]), .IN2(n43), .IN3(data0[9]), .IN4(n42), .IN5(n41), 
        .Q(data_o[9]) );
  AO22X1 U6 ( .IN1(data2[9]), .IN2(n40), .IN3(data3[9]), .IN4(n39), .Q(n41) );
  AO221X1 U7 ( .IN1(data1[8]), .IN2(n43), .IN3(data0[8]), .IN4(n42), .IN5(n38), 
        .Q(data_o[8]) );
  AO22X1 U8 ( .IN1(data2[8]), .IN2(n40), .IN3(data3[8]), .IN4(n39), .Q(n38) );
  AO221X1 U9 ( .IN1(data1[7]), .IN2(n43), .IN3(data0[7]), .IN4(n42), .IN5(n37), 
        .Q(data_o[7]) );
  AO22X1 U10 ( .IN1(data2[7]), .IN2(n40), .IN3(data3[7]), .IN4(n39), .Q(n37)
         );
  AO221X1 U11 ( .IN1(data1[6]), .IN2(n43), .IN3(data0[6]), .IN4(n42), .IN5(n36), .Q(data_o[6]) );
  AO22X1 U12 ( .IN1(data2[6]), .IN2(n40), .IN3(data3[6]), .IN4(n39), .Q(n36)
         );
  AO221X1 U13 ( .IN1(data1[5]), .IN2(n43), .IN3(data0[5]), .IN4(n42), .IN5(n35), .Q(data_o[5]) );
  AO22X1 U14 ( .IN1(data2[5]), .IN2(n40), .IN3(data3[5]), .IN4(n39), .Q(n35)
         );
  AO221X1 U15 ( .IN1(data1[4]), .IN2(n43), .IN3(data0[4]), .IN4(n42), .IN5(n34), .Q(data_o[4]) );
  AO22X1 U16 ( .IN1(data2[4]), .IN2(n40), .IN3(data3[4]), .IN4(n39), .Q(n34)
         );
  AO221X1 U17 ( .IN1(data1[3]), .IN2(n43), .IN3(data0[3]), .IN4(n42), .IN5(n33), .Q(data_o[3]) );
  AO22X1 U18 ( .IN1(data2[3]), .IN2(n40), .IN3(data3[3]), .IN4(n39), .Q(n33)
         );
  AO221X1 U19 ( .IN1(data1[2]), .IN2(n43), .IN3(data0[2]), .IN4(n42), .IN5(n32), .Q(data_o[2]) );
  AO22X1 U20 ( .IN1(data2[2]), .IN2(n40), .IN3(data3[2]), .IN4(n39), .Q(n32)
         );
  AO221X1 U21 ( .IN1(data1[1]), .IN2(n43), .IN3(data0[1]), .IN4(n42), .IN5(n31), .Q(data_o[1]) );
  AO22X1 U22 ( .IN1(data2[1]), .IN2(n40), .IN3(data3[1]), .IN4(n39), .Q(n31)
         );
  AO221X1 U23 ( .IN1(data1[15]), .IN2(n43), .IN3(data0[15]), .IN4(n42), .IN5(
        n30), .Q(data_o[15]) );
  AO22X1 U24 ( .IN1(data2[15]), .IN2(n40), .IN3(data3[15]), .IN4(n39), .Q(n30)
         );
  AO221X1 U25 ( .IN1(data1[14]), .IN2(n43), .IN3(data0[14]), .IN4(n42), .IN5(
        n29), .Q(data_o[14]) );
  AO22X1 U26 ( .IN1(data2[14]), .IN2(n40), .IN3(data3[14]), .IN4(n39), .Q(n29)
         );
  AO221X1 U27 ( .IN1(data1[13]), .IN2(n43), .IN3(data0[13]), .IN4(n42), .IN5(
        n28), .Q(data_o[13]) );
  AO22X1 U28 ( .IN1(data2[13]), .IN2(n40), .IN3(data3[13]), .IN4(n39), .Q(n28)
         );
  AO221X1 U29 ( .IN1(data1[12]), .IN2(n43), .IN3(data0[12]), .IN4(n42), .IN5(
        n27), .Q(data_o[12]) );
  AO22X1 U30 ( .IN1(data2[12]), .IN2(n40), .IN3(data3[12]), .IN4(n39), .Q(n27)
         );
  AO221X1 U31 ( .IN1(data1[11]), .IN2(n43), .IN3(data0[11]), .IN4(n42), .IN5(
        n26), .Q(data_o[11]) );
  AO22X1 U32 ( .IN1(data2[11]), .IN2(n40), .IN3(data3[11]), .IN4(n39), .Q(n26)
         );
  AO221X1 U33 ( .IN1(data1[10]), .IN2(n43), .IN3(data0[10]), .IN4(n42), .IN5(
        n25), .Q(data_o[10]) );
  AO22X1 U34 ( .IN1(data2[10]), .IN2(n40), .IN3(data3[10]), .IN4(n39), .Q(n25)
         );
  AO221X1 U35 ( .IN1(data1[0]), .IN2(n43), .IN3(data0[0]), .IN4(n42), .IN5(n24), .Q(data_o[0]) );
  AO22X1 U36 ( .IN1(data2[0]), .IN2(n40), .IN3(data3[0]), .IN4(n39), .Q(n24)
         );
  INVX0 U2 ( .INP(select2), .ZN(n1) );
  NOR4X0 U3 ( .IN1(n1), .IN2(select0), .IN3(select1), .IN4(select3), .QN(n40)
         );
  AND4X1 U4 ( .IN1(select3), .IN2(n3), .IN3(n2), .IN4(n1), .Q(n39) );
  INVX0 U37 ( .INP(select0), .ZN(n3) );
  INVX0 U38 ( .INP(select1), .ZN(n2) );
  NOR4X0 U39 ( .IN1(n3), .IN2(select1), .IN3(select2), .IN4(select3), .QN(n42)
         );
  NOR4X0 U40 ( .IN1(n2), .IN2(select0), .IN3(select2), .IN4(select3), .QN(n43)
         );
endmodule


module mux4_1_0 ( data0, data1, data2, data3, select0, select1, select2, 
        select3, data_o );
  input [15:0] data0;
  input [15:0] data1;
  input [15:0] data2;
  input [15:0] data3;
  output [15:0] data_o;
  input select0, select1, select2, select3;
  wire   n1, n2, n3, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43;

  AO221X1 U5 ( .IN1(data1[9]), .IN2(n43), .IN3(data0[9]), .IN4(n42), .IN5(n41), 
        .Q(data_o[9]) );
  AO22X1 U6 ( .IN1(data2[9]), .IN2(n40), .IN3(data3[9]), .IN4(n39), .Q(n41) );
  AO221X1 U7 ( .IN1(data1[8]), .IN2(n43), .IN3(data0[8]), .IN4(n42), .IN5(n38), 
        .Q(data_o[8]) );
  AO22X1 U8 ( .IN1(data2[8]), .IN2(n40), .IN3(data3[8]), .IN4(n39), .Q(n38) );
  AO221X1 U9 ( .IN1(data1[7]), .IN2(n43), .IN3(data0[7]), .IN4(n42), .IN5(n37), 
        .Q(data_o[7]) );
  AO22X1 U10 ( .IN1(data2[7]), .IN2(n40), .IN3(data3[7]), .IN4(n39), .Q(n37)
         );
  AO221X1 U11 ( .IN1(data1[6]), .IN2(n43), .IN3(data0[6]), .IN4(n42), .IN5(n36), .Q(data_o[6]) );
  AO22X1 U12 ( .IN1(data2[6]), .IN2(n40), .IN3(data3[6]), .IN4(n39), .Q(n36)
         );
  AO221X1 U13 ( .IN1(data1[5]), .IN2(n43), .IN3(data0[5]), .IN4(n42), .IN5(n35), .Q(data_o[5]) );
  AO22X1 U14 ( .IN1(data2[5]), .IN2(n40), .IN3(data3[5]), .IN4(n39), .Q(n35)
         );
  AO221X1 U15 ( .IN1(data1[4]), .IN2(n43), .IN3(data0[4]), .IN4(n42), .IN5(n34), .Q(data_o[4]) );
  AO22X1 U16 ( .IN1(data2[4]), .IN2(n40), .IN3(data3[4]), .IN4(n39), .Q(n34)
         );
  AO221X1 U17 ( .IN1(data1[3]), .IN2(n43), .IN3(data0[3]), .IN4(n42), .IN5(n33), .Q(data_o[3]) );
  AO22X1 U18 ( .IN1(data2[3]), .IN2(n40), .IN3(data3[3]), .IN4(n39), .Q(n33)
         );
  AO221X1 U19 ( .IN1(data1[2]), .IN2(n43), .IN3(data0[2]), .IN4(n42), .IN5(n32), .Q(data_o[2]) );
  AO22X1 U20 ( .IN1(data2[2]), .IN2(n40), .IN3(data3[2]), .IN4(n39), .Q(n32)
         );
  AO221X1 U21 ( .IN1(data1[1]), .IN2(n43), .IN3(data0[1]), .IN4(n42), .IN5(n31), .Q(data_o[1]) );
  AO22X1 U22 ( .IN1(data2[1]), .IN2(n40), .IN3(data3[1]), .IN4(n39), .Q(n31)
         );
  AO221X1 U23 ( .IN1(data1[15]), .IN2(n43), .IN3(data0[15]), .IN4(n42), .IN5(
        n30), .Q(data_o[15]) );
  AO22X1 U24 ( .IN1(data2[15]), .IN2(n40), .IN3(data3[15]), .IN4(n39), .Q(n30)
         );
  AO221X1 U25 ( .IN1(data1[14]), .IN2(n43), .IN3(data0[14]), .IN4(n42), .IN5(
        n29), .Q(data_o[14]) );
  AO22X1 U26 ( .IN1(data2[14]), .IN2(n40), .IN3(data3[14]), .IN4(n39), .Q(n29)
         );
  AO221X1 U27 ( .IN1(data1[13]), .IN2(n43), .IN3(data0[13]), .IN4(n42), .IN5(
        n28), .Q(data_o[13]) );
  AO22X1 U28 ( .IN1(data2[13]), .IN2(n40), .IN3(data3[13]), .IN4(n39), .Q(n28)
         );
  AO221X1 U29 ( .IN1(data1[12]), .IN2(n43), .IN3(data0[12]), .IN4(n42), .IN5(
        n27), .Q(data_o[12]) );
  AO22X1 U30 ( .IN1(data2[12]), .IN2(n40), .IN3(data3[12]), .IN4(n39), .Q(n27)
         );
  AO221X1 U31 ( .IN1(data1[11]), .IN2(n43), .IN3(data0[11]), .IN4(n42), .IN5(
        n26), .Q(data_o[11]) );
  AO22X1 U32 ( .IN1(data2[11]), .IN2(n40), .IN3(data3[11]), .IN4(n39), .Q(n26)
         );
  AO221X1 U33 ( .IN1(data1[10]), .IN2(n43), .IN3(data0[10]), .IN4(n42), .IN5(
        n25), .Q(data_o[10]) );
  AO22X1 U34 ( .IN1(data2[10]), .IN2(n40), .IN3(data3[10]), .IN4(n39), .Q(n25)
         );
  AO221X1 U35 ( .IN1(data1[0]), .IN2(n43), .IN3(data0[0]), .IN4(n42), .IN5(n24), .Q(data_o[0]) );
  AO22X1 U36 ( .IN1(data2[0]), .IN2(n40), .IN3(data3[0]), .IN4(n39), .Q(n24)
         );
  INVX0 U2 ( .INP(select2), .ZN(n1) );
  NOR4X0 U3 ( .IN1(n1), .IN2(select0), .IN3(select1), .IN4(select3), .QN(n40)
         );
  AND4X1 U4 ( .IN1(select3), .IN2(n3), .IN3(n2), .IN4(n1), .Q(n39) );
  INVX0 U37 ( .INP(select0), .ZN(n3) );
  INVX0 U38 ( .INP(select1), .ZN(n2) );
  NOR4X0 U39 ( .IN1(n3), .IN2(select1), .IN3(select2), .IN4(select3), .QN(n42)
         );
  NOR4X0 U40 ( .IN1(n2), .IN2(select0), .IN3(select2), .IN4(select3), .QN(n43)
         );
endmodule



    module node5_NODE_X2_NODE_Y2I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__I_node_2_node_interface__I_node_3_node_interface__ ( 
        \clk.clk , \reset.reset , \local_node.clk , 
        \local_node.buffer_full_in , \local_node.buffer_full_out , 
        \local_node.receiving_data , \local_node.sending_data , 
        \local_node.data_in , \local_node.data_out , \node_0.clk , 
        \node_0.buffer_full_in , \node_0.buffer_full_out , 
        \node_0.receiving_data , \node_0.sending_data , \node_0.data_in , 
        \node_0.data_out , \node_1.clk , \node_1.buffer_full_in , 
        \node_1.buffer_full_out , \node_1.receiving_data , 
        \node_1.sending_data , \node_1.data_in , \node_1.data_out , 
        \node_2.clk , \node_2.buffer_full_in , \node_2.buffer_full_out , 
        \node_2.receiving_data , \node_2.sending_data , \node_2.data_in , 
        \node_2.data_out , \node_3.clk , \node_3.buffer_full_in , 
        \node_3.buffer_full_out , \node_3.receiving_data , 
        \node_3.sending_data , \node_3.data_in , \node_3.data_out  );
  input [15:0] \local_node.data_in ;
  output [15:0] \local_node.data_out ;
  input [15:0] \node_0.data_in ;
  output [15:0] \node_0.data_out ;
  input [15:0] \node_1.data_in ;
  output [15:0] \node_1.data_out ;
  input [15:0] \node_2.data_in ;
  output [15:0] \node_2.data_out ;
  input [15:0] \node_3.data_in ;
  output [15:0] \node_3.data_out ;
  input \clk.clk , \reset.reset , \local_node.buffer_full_in ,
         \local_node.receiving_data , \node_0.buffer_full_in ,
         \node_0.receiving_data , \node_1.buffer_full_in ,
         \node_1.receiving_data , \node_2.buffer_full_in ,
         \node_2.receiving_data , \node_3.buffer_full_in ,
         \node_3.receiving_data ;
  output \local_node.buffer_full_out , \local_node.sending_data ,
         \node_0.buffer_full_out , \node_0.sending_data ,
         \node_1.buffer_full_out , \node_1.sending_data ,
         \node_2.buffer_full_out , \node_2.sending_data ,
         \node_3.buffer_full_out , \node_3.sending_data ;
  inout \local_node.clk ,  \node_0.clk ,  \node_1.clk ,  \node_2.clk , 
     \node_3.clk ;
  wire   \buffer_out[4][15] , \buffer_out[4][14] , \buffer_out[4][13] ,
         \buffer_out[4][12] , \buffer_out[4][11] , \buffer_out[4][10] ,
         \buffer_out[4][9] , \buffer_out[4][8] , \buffer_out[4][7] ,
         \buffer_out[4][6] , \buffer_out[4][5] , \buffer_out[4][4] ,
         \buffer_out[4][3] , \buffer_out[4][2] , \buffer_out[4][1] ,
         \buffer_out[4][0] , \buffer_out[3][15] , \buffer_out[3][14] ,
         \buffer_out[3][13] , \buffer_out[3][12] , \buffer_out[3][11] ,
         \buffer_out[3][10] , \buffer_out[3][9] , \buffer_out[3][8] ,
         \buffer_out[3][7] , \buffer_out[3][6] , \buffer_out[3][5] ,
         \buffer_out[3][4] , \buffer_out[3][3] , \buffer_out[3][2] ,
         \buffer_out[3][1] , \buffer_out[3][0] , \buffer_out[2][15] ,
         \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] ,
         \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] ,
         \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] ,
         \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] ,
         \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] ,
         \buffer_out[1][15] , \buffer_out[1][14] , \buffer_out[1][13] ,
         \buffer_out[1][12] , \buffer_out[1][11] , \buffer_out[1][10] ,
         \buffer_out[1][9] , \buffer_out[1][8] , \buffer_out[1][7] ,
         \buffer_out[1][6] , \buffer_out[1][5] , \buffer_out[1][4] ,
         \buffer_out[1][3] , \buffer_out[1][2] , \buffer_out[1][1] ,
         \buffer_out[1][0] , \buffer_out[0][15] , \buffer_out[0][14] ,
         \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] ,
         \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] ,
         \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] ,
         \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] ,
         \buffer_out[0][1] , \buffer_out[0][0] , \next_buffer_out[4][15] ,
         \next_buffer_out[4][14] , \next_buffer_out[4][13] ,
         \next_buffer_out[4][12] , \next_buffer_out[4][11] ,
         \next_buffer_out[4][10] , \next_buffer_out[4][9] ,
         \next_buffer_out[4][8] , \next_buffer_out[4][7] ,
         \next_buffer_out[4][6] , \next_buffer_out[4][5] ,
         \next_buffer_out[4][4] , \next_buffer_out[4][3] ,
         \next_buffer_out[4][2] , \next_buffer_out[4][1] ,
         \next_buffer_out[4][0] , \next_buffer_out[3][15] ,
         \next_buffer_out[3][14] , \next_buffer_out[3][13] ,
         \next_buffer_out[3][12] , \next_buffer_out[3][11] ,
         \next_buffer_out[3][10] , \next_buffer_out[3][9] ,
         \next_buffer_out[3][8] , \next_buffer_out[3][7] ,
         \next_buffer_out[3][6] , \next_buffer_out[3][5] ,
         \next_buffer_out[3][4] , \next_buffer_out[3][3] ,
         \next_buffer_out[3][2] , \next_buffer_out[3][1] ,
         \next_buffer_out[3][0] , \next_buffer_out[2][15] ,
         \next_buffer_out[2][14] , \next_buffer_out[2][13] ,
         \next_buffer_out[2][12] , \next_buffer_out[2][11] ,
         \next_buffer_out[2][10] , \next_buffer_out[2][9] ,
         \next_buffer_out[2][8] , \next_buffer_out[2][7] ,
         \next_buffer_out[2][6] , \next_buffer_out[2][5] ,
         \next_buffer_out[2][4] , \next_buffer_out[2][3] ,
         \next_buffer_out[2][2] , \next_buffer_out[2][1] ,
         \next_buffer_out[2][0] , \next_buffer_out[1][15] ,
         \next_buffer_out[1][14] , \next_buffer_out[1][13] ,
         \next_buffer_out[1][12] , \next_buffer_out[1][11] ,
         \next_buffer_out[1][10] , \next_buffer_out[1][9] ,
         \next_buffer_out[1][8] , \next_buffer_out[1][7] ,
         \next_buffer_out[1][6] , \next_buffer_out[1][5] ,
         \next_buffer_out[1][4] , \next_buffer_out[1][3] ,
         \next_buffer_out[1][2] , \next_buffer_out[1][1] ,
         \next_buffer_out[1][0] , \next_buffer_out[0][15] ,
         \next_buffer_out[0][14] , \next_buffer_out[0][13] ,
         \next_buffer_out[0][12] , \next_buffer_out[0][11] ,
         \next_buffer_out[0][10] , \next_buffer_out[0][9] ,
         \next_buffer_out[0][8] , \next_buffer_out[0][7] ,
         \next_buffer_out[0][6] , \next_buffer_out[0][5] ,
         \next_buffer_out[0][4] , \next_buffer_out[0][3] ,
         \next_buffer_out[0][2] , \next_buffer_out[0][1] ,
         \next_buffer_out[0][0] ;
  wire   [4:0] buffer_full_in;
  wire   [4:0] receiving_data;
  wire   [4:0] pop_v;
  wire   [4:0] data_valid;
  wire   [4:0] next_data_valid;
  wire   [1:0] grant_0;
  wire   [1:0] grant_1;
  wire   [3:0] grant_2;
  wire   [3:0] grant_3;
  wire   [3:0] grant_4;
  tri   \local_node.buffer_full_in ;
  tri   \local_node.buffer_full_out ;
  tri   \local_node.receiving_data ;
  tri   \local_node.sending_data ;
  tri   [15:0] \local_node.data_in ;
  tri   [15:0] \local_node.data_out ;

  converter_in_I_n_node_interface_dut__1 c0 ( .\n.buffer_full_in (
        \node_0.buffer_full_in ), .\n.receiving_data (\node_0.receiving_data ), 
        .\n.data_in (\node_0.data_in ), .\n.buffer_full_out (
        \node_0.buffer_full_out ), .\n.sending_data (\node_0.sending_data ), 
        .\n.data_out (\node_0.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_out_I_n_node_interface_dut_ c1 ( .\n.buffer_full_in (
        \node_1.buffer_full_in ), .\n.receiving_data (\node_1.receiving_data ), 
        .\n.data_in (\node_1.data_in ), .\n.buffer_full_out (
        \node_1.buffer_full_out ), .\n.sending_data (\node_1.sending_data ), 
        .\n.data_out (\node_1.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_in_I_n_node_interface_dut__0 c2 ( .\n.buffer_full_in (
        \node_2.buffer_full_in ), .\n.receiving_data (\node_2.receiving_data ), 
        .\n.data_in (\node_2.data_in ), .\n.buffer_full_out (
        \node_2.buffer_full_out ), .\n.sending_data (\node_2.sending_data ), 
        .\n.data_out (\node_2.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_out_I_n_node_interface_dut_ c3 ( .\n.buffer_full_in (
        \node_3.buffer_full_in ), .\n.receiving_data (\node_3.receiving_data ), 
        .\n.data_in (\node_3.data_in ), .\n.buffer_full_out (
        \node_3.buffer_full_out ), .\n.sending_data (\node_3.sending_data ), 
        .\n.data_out (\node_3.data_out ), .buffer_full_in(1'b0), 
        .receiving_data(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  converter_out_I_n_node_interface_dut_ c4 ( .\n.buffer_full_in (
        \local_node.buffer_full_in ), .\n.receiving_data (
        \local_node.receiving_data ), .\n.data_in (\local_node.data_in ), 
        .\n.buffer_full_out (\local_node.buffer_full_out ), .\n.sending_data (
        \local_node.sending_data ), .\n.data_out (\local_node.data_out ), 
        .buffer_full_in(1'b0), .receiving_data(1'b0), .data_in({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  fifo_kev_4 \genblk1[0].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[0]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[0]), .data_out({\buffer_out[0][15] , 
        \buffer_out[0][14] , \buffer_out[0][13] , \buffer_out[0][12] , 
        \buffer_out[0][11] , \buffer_out[0][10] , \buffer_out[0][9] , 
        \buffer_out[0][8] , \buffer_out[0][7] , \buffer_out[0][6] , 
        \buffer_out[0][5] , \buffer_out[0][4] , \buffer_out[0][3] , 
        \buffer_out[0][2] , \buffer_out[0][1] , \buffer_out[0][0] }), 
        .next_data_out({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] , 
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .next_data_valid(
        next_data_valid[0]) );
  address_counter_4 \genblk1[0].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[0][15] , \next_buffer_out[0][14] , 
        \next_buffer_out[0][13] , \next_buffer_out[0][12] , 
        \next_buffer_out[0][11] , \next_buffer_out[0][10] , 
        \next_buffer_out[0][9] , \next_buffer_out[0][8] }), 
        .buffer_data_valid(next_data_valid[0]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[0][7] , \next_buffer_out[0][6] , 
        \next_buffer_out[0][5] , \next_buffer_out[0][4] , 
        \next_buffer_out[0][3] , \next_buffer_out[0][2] , 
        \next_buffer_out[0][1] , \next_buffer_out[0][0] }), .buffer_pop(
        pop_v[0]), .receiving_data(1'b0) );
  fifo_kev_3 \genblk1[1].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[1]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[1]), .data_out({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), 
        .next_data_out({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] , 
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .next_data_valid(
        next_data_valid[1]) );
  address_counter_3 \genblk1[1].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[1][15] , \next_buffer_out[1][14] , 
        \next_buffer_out[1][13] , \next_buffer_out[1][12] , 
        \next_buffer_out[1][11] , \next_buffer_out[1][10] , 
        \next_buffer_out[1][9] , \next_buffer_out[1][8] }), 
        .buffer_data_valid(next_data_valid[1]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[1][7] , \next_buffer_out[1][6] , 
        \next_buffer_out[1][5] , \next_buffer_out[1][4] , 
        \next_buffer_out[1][3] , \next_buffer_out[1][2] , 
        \next_buffer_out[1][1] , \next_buffer_out[1][0] }), .buffer_pop(
        pop_v[1]), .receiving_data(1'b0) );
  fifo_kev_2 \genblk1[2].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[2]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[2]), .data_out({\buffer_out[2][15] , 
        \buffer_out[2][14] , \buffer_out[2][13] , \buffer_out[2][12] , 
        \buffer_out[2][11] , \buffer_out[2][10] , \buffer_out[2][9] , 
        \buffer_out[2][8] , \buffer_out[2][7] , \buffer_out[2][6] , 
        \buffer_out[2][5] , \buffer_out[2][4] , \buffer_out[2][3] , 
        \buffer_out[2][2] , \buffer_out[2][1] , \buffer_out[2][0] }), 
        .next_data_out({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] , 
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .next_data_valid(
        next_data_valid[2]) );
  address_counter_2 \genblk1[2].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[2][15] , \next_buffer_out[2][14] , 
        \next_buffer_out[2][13] , \next_buffer_out[2][12] , 
        \next_buffer_out[2][11] , \next_buffer_out[2][10] , 
        \next_buffer_out[2][9] , \next_buffer_out[2][8] }), 
        .buffer_data_valid(next_data_valid[2]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[2][7] , \next_buffer_out[2][6] , 
        \next_buffer_out[2][5] , \next_buffer_out[2][4] , 
        \next_buffer_out[2][3] , \next_buffer_out[2][2] , 
        \next_buffer_out[2][1] , \next_buffer_out[2][0] }), .buffer_pop(
        pop_v[2]), .receiving_data(1'b0) );
  fifo_kev_1 \genblk1[3].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[3]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[3]), .data_out({\buffer_out[3][15] , 
        \buffer_out[3][14] , \buffer_out[3][13] , \buffer_out[3][12] , 
        \buffer_out[3][11] , \buffer_out[3][10] , \buffer_out[3][9] , 
        \buffer_out[3][8] , \buffer_out[3][7] , \buffer_out[3][6] , 
        \buffer_out[3][5] , \buffer_out[3][4] , \buffer_out[3][3] , 
        \buffer_out[3][2] , \buffer_out[3][1] , \buffer_out[3][0] }), 
        .next_data_out({\next_buffer_out[3][15] , \next_buffer_out[3][14] , 
        \next_buffer_out[3][13] , \next_buffer_out[3][12] , 
        \next_buffer_out[3][11] , \next_buffer_out[3][10] , 
        \next_buffer_out[3][9] , \next_buffer_out[3][8] , 
        \next_buffer_out[3][7] , \next_buffer_out[3][6] , 
        \next_buffer_out[3][5] , \next_buffer_out[3][4] , 
        \next_buffer_out[3][3] , \next_buffer_out[3][2] , 
        \next_buffer_out[3][1] , \next_buffer_out[3][0] }), .next_data_valid(
        next_data_valid[3]) );
  address_counter_1 \genblk1[3].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[3][15] , \next_buffer_out[3][14] , 
        \next_buffer_out[3][13] , \next_buffer_out[3][12] , 
        \next_buffer_out[3][11] , \next_buffer_out[3][10] , 
        \next_buffer_out[3][9] , \next_buffer_out[3][8] }), 
        .buffer_data_valid(next_data_valid[3]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[3][7] , \next_buffer_out[3][6] , 
        \next_buffer_out[3][5] , \next_buffer_out[3][4] , 
        \next_buffer_out[3][3] , \next_buffer_out[3][2] , 
        \next_buffer_out[3][1] , \next_buffer_out[3][0] }), .buffer_pop(
        pop_v[3]), .receiving_data(1'b0) );
  fifo_kev_0 \genblk1[4].buffer  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .push_req(1'b0), .pop_req(pop_v[4]), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .data_valid(data_valid[4]), .data_out({\buffer_out[4][15] , 
        \buffer_out[4][14] , \buffer_out[4][13] , \buffer_out[4][12] , 
        \buffer_out[4][11] , \buffer_out[4][10] , \buffer_out[4][9] , 
        \buffer_out[4][8] , \buffer_out[4][7] , \buffer_out[4][6] , 
        \buffer_out[4][5] , \buffer_out[4][4] , \buffer_out[4][3] , 
        \buffer_out[4][2] , \buffer_out[4][1] , \buffer_out[4][0] }), 
        .next_data_out({\next_buffer_out[4][15] , \next_buffer_out[4][14] , 
        \next_buffer_out[4][13] , \next_buffer_out[4][12] , 
        \next_buffer_out[4][11] , \next_buffer_out[4][10] , 
        \next_buffer_out[4][9] , \next_buffer_out[4][8] , 
        \next_buffer_out[4][7] , \next_buffer_out[4][6] , 
        \next_buffer_out[4][5] , \next_buffer_out[4][4] , 
        \next_buffer_out[4][3] , \next_buffer_out[4][2] , 
        \next_buffer_out[4][1] , \next_buffer_out[4][0] }), .next_data_valid(
        next_data_valid[4]) );
  address_counter_0 \genblk1[4].addr  ( .clk(\clk.clk ), .rst(\reset.reset ), 
        .interface_flit_length({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_length({\next_buffer_out[4][15] , \next_buffer_out[4][14] , 
        \next_buffer_out[4][13] , \next_buffer_out[4][12] , 
        \next_buffer_out[4][11] , \next_buffer_out[4][10] , 
        \next_buffer_out[4][9] , \next_buffer_out[4][8] }), 
        .buffer_data_valid(next_data_valid[4]), .interface_flit_address({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .buffer_flit_address({
        \next_buffer_out[4][7] , \next_buffer_out[4][6] , 
        \next_buffer_out[4][5] , \next_buffer_out[4][4] , 
        \next_buffer_out[4][3] , \next_buffer_out[4][2] , 
        \next_buffer_out[4][1] , \next_buffer_out[4][0] }), .buffer_pop(
        pop_v[4]), .receiving_data(1'b0) );
  controller5_0 ctrl5 ( .clk(\clk.clk ), .rst(\reset.reset ), .packet_addr({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .local_addr({1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 
        1'b0, 1'b1, 1'b0}), .packet_valid(data_valid), .buffer_full_in({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .grant_0(grant_0), .grant_1(grant_1), 
        .grant_2(grant_2), .grant_3(grant_3), .grant_4(grant_4), .pop_v(pop_v)
         );
  mux2_1_1 mux_n ( .data0({\buffer_out[1][15] , \buffer_out[1][14] , 
        \buffer_out[1][13] , \buffer_out[1][12] , \buffer_out[1][11] , 
        \buffer_out[1][10] , \buffer_out[1][9] , \buffer_out[1][8] , 
        \buffer_out[1][7] , \buffer_out[1][6] , \buffer_out[1][5] , 
        \buffer_out[1][4] , \buffer_out[1][3] , \buffer_out[1][2] , 
        \buffer_out[1][1] , \buffer_out[1][0] }), .data1({\buffer_out[4][15] , 
        \buffer_out[4][14] , \buffer_out[4][13] , \buffer_out[4][12] , 
        \buffer_out[4][11] , \buffer_out[4][10] , \buffer_out[4][9] , 
        \buffer_out[4][8] , \buffer_out[4][7] , \buffer_out[4][6] , 
        \buffer_out[4][5] , \buffer_out[4][4] , \buffer_out[4][3] , 
        \buffer_out[4][2] , \buffer_out[4][1] , \buffer_out[4][0] }), 
        .select0(grant_0[0]), .select1(grant_0[1]) );
  mux2_1_0 mux_s ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[4][15] , 
        \buffer_out[4][14] , \buffer_out[4][13] , \buffer_out[4][12] , 
        \buffer_out[4][11] , \buffer_out[4][10] , \buffer_out[4][9] , 
        \buffer_out[4][8] , \buffer_out[4][7] , \buffer_out[4][6] , 
        \buffer_out[4][5] , \buffer_out[4][4] , \buffer_out[4][3] , 
        \buffer_out[4][2] , \buffer_out[4][1] , \buffer_out[4][0] }), 
        .select0(grant_1[0]), .select1(grant_1[1]) );
  mux4_1_2 mux_e ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[3][15] , \buffer_out[3][14] , \buffer_out[3][13] , 
        \buffer_out[3][12] , \buffer_out[3][11] , \buffer_out[3][10] , 
        \buffer_out[3][9] , \buffer_out[3][8] , \buffer_out[3][7] , 
        \buffer_out[3][6] , \buffer_out[3][5] , \buffer_out[3][4] , 
        \buffer_out[3][3] , \buffer_out[3][2] , \buffer_out[3][1] , 
        \buffer_out[3][0] }), .data3({\buffer_out[4][15] , \buffer_out[4][14] , 
        \buffer_out[4][13] , \buffer_out[4][12] , \buffer_out[4][11] , 
        \buffer_out[4][10] , \buffer_out[4][9] , \buffer_out[4][8] , 
        \buffer_out[4][7] , \buffer_out[4][6] , \buffer_out[4][5] , 
        \buffer_out[4][4] , \buffer_out[4][3] , \buffer_out[4][2] , 
        \buffer_out[4][1] , \buffer_out[4][0] }), .select0(grant_2[0]), 
        .select1(grant_2[1]), .select2(grant_2[2]), .select3(grant_2[3]) );
  mux4_1_1 mux_w ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[2][15] , \buffer_out[2][14] , \buffer_out[2][13] , 
        \buffer_out[2][12] , \buffer_out[2][11] , \buffer_out[2][10] , 
        \buffer_out[2][9] , \buffer_out[2][8] , \buffer_out[2][7] , 
        \buffer_out[2][6] , \buffer_out[2][5] , \buffer_out[2][4] , 
        \buffer_out[2][3] , \buffer_out[2][2] , \buffer_out[2][1] , 
        \buffer_out[2][0] }), .data3({\buffer_out[4][15] , \buffer_out[4][14] , 
        \buffer_out[4][13] , \buffer_out[4][12] , \buffer_out[4][11] , 
        \buffer_out[4][10] , \buffer_out[4][9] , \buffer_out[4][8] , 
        \buffer_out[4][7] , \buffer_out[4][6] , \buffer_out[4][5] , 
        \buffer_out[4][4] , \buffer_out[4][3] , \buffer_out[4][2] , 
        \buffer_out[4][1] , \buffer_out[4][0] }), .select0(grant_3[0]), 
        .select1(grant_3[1]), .select2(grant_3[2]), .select3(grant_3[3]) );
  mux4_1_0 mux_l ( .data0({\buffer_out[0][15] , \buffer_out[0][14] , 
        \buffer_out[0][13] , \buffer_out[0][12] , \buffer_out[0][11] , 
        \buffer_out[0][10] , \buffer_out[0][9] , \buffer_out[0][8] , 
        \buffer_out[0][7] , \buffer_out[0][6] , \buffer_out[0][5] , 
        \buffer_out[0][4] , \buffer_out[0][3] , \buffer_out[0][2] , 
        \buffer_out[0][1] , \buffer_out[0][0] }), .data1({\buffer_out[1][15] , 
        \buffer_out[1][14] , \buffer_out[1][13] , \buffer_out[1][12] , 
        \buffer_out[1][11] , \buffer_out[1][10] , \buffer_out[1][9] , 
        \buffer_out[1][8] , \buffer_out[1][7] , \buffer_out[1][6] , 
        \buffer_out[1][5] , \buffer_out[1][4] , \buffer_out[1][3] , 
        \buffer_out[1][2] , \buffer_out[1][1] , \buffer_out[1][0] }), .data2({
        \buffer_out[2][15] , \buffer_out[2][14] , \buffer_out[2][13] , 
        \buffer_out[2][12] , \buffer_out[2][11] , \buffer_out[2][10] , 
        \buffer_out[2][9] , \buffer_out[2][8] , \buffer_out[2][7] , 
        \buffer_out[2][6] , \buffer_out[2][5] , \buffer_out[2][4] , 
        \buffer_out[2][3] , \buffer_out[2][2] , \buffer_out[2][1] , 
        \buffer_out[2][0] }), .data3({\buffer_out[3][15] , \buffer_out[3][14] , 
        \buffer_out[3][13] , \buffer_out[3][12] , \buffer_out[3][11] , 
        \buffer_out[3][10] , \buffer_out[3][9] , \buffer_out[3][8] , 
        \buffer_out[3][7] , \buffer_out[3][6] , \buffer_out[3][5] , 
        \buffer_out[3][4] , \buffer_out[3][3] , \buffer_out[3][2] , 
        \buffer_out[3][1] , \buffer_out[3][0] }), .select0(grant_4[0]), 
        .select1(grant_4[1]), .select2(grant_4[2]), .select3(grant_4[3]) );
endmodule


module noc ( \clk.clk , \reset.reset , \local_node[0].clk , 
        \local_node[0].buffer_full_in , \local_node[0].buffer_full_out , 
        \local_node[0].receiving_data , \local_node[0].sending_data , 
        \local_node[0].data_in , \local_node[0].data_out , \local_node[1].clk , 
        \local_node[1].buffer_full_in , \local_node[1].buffer_full_out , 
        \local_node[1].receiving_data , \local_node[1].sending_data , 
        \local_node[1].data_in , \local_node[1].data_out , \local_node[2].clk , 
        \local_node[2].buffer_full_in , \local_node[2].buffer_full_out , 
        \local_node[2].receiving_data , \local_node[2].sending_data , 
        \local_node[2].data_in , \local_node[2].data_out , \local_node[3].clk , 
        \local_node[3].buffer_full_in , \local_node[3].buffer_full_out , 
        \local_node[3].receiving_data , \local_node[3].sending_data , 
        \local_node[3].data_in , \local_node[3].data_out , \local_node[4].clk , 
        \local_node[4].buffer_full_in , \local_node[4].buffer_full_out , 
        \local_node[4].receiving_data , \local_node[4].sending_data , 
        \local_node[4].data_in , \local_node[4].data_out , \local_node[5].clk , 
        \local_node[5].buffer_full_in , \local_node[5].buffer_full_out , 
        \local_node[5].receiving_data , \local_node[5].sending_data , 
        \local_node[5].data_in , \local_node[5].data_out , \local_node[6].clk , 
        \local_node[6].buffer_full_in , \local_node[6].buffer_full_out , 
        \local_node[6].receiving_data , \local_node[6].sending_data , 
        \local_node[6].data_in , \local_node[6].data_out , \local_node[7].clk , 
        \local_node[7].buffer_full_in , \local_node[7].buffer_full_out , 
        \local_node[7].receiving_data , \local_node[7].sending_data , 
        \local_node[7].data_in , \local_node[7].data_out , \local_node[8].clk , 
        \local_node[8].buffer_full_in , \local_node[8].buffer_full_out , 
        \local_node[8].receiving_data , \local_node[8].sending_data , 
        \local_node[8].data_in , \local_node[8].data_out , \local_node[9].clk , 
        \local_node[9].buffer_full_in , \local_node[9].buffer_full_out , 
        \local_node[9].receiving_data , \local_node[9].sending_data , 
        \local_node[9].data_in , \local_node[9].data_out , 
        \local_node[10].clk , \local_node[10].buffer_full_in , 
        \local_node[10].buffer_full_out , \local_node[10].receiving_data , 
        \local_node[10].sending_data , \local_node[10].data_in , 
        \local_node[10].data_out , \local_node[11].clk , 
        \local_node[11].buffer_full_in , \local_node[11].buffer_full_out , 
        \local_node[11].receiving_data , \local_node[11].sending_data , 
        \local_node[11].data_in , \local_node[11].data_out , 
        \local_node[12].clk , \local_node[12].buffer_full_in , 
        \local_node[12].buffer_full_out , \local_node[12].receiving_data , 
        \local_node[12].sending_data , \local_node[12].data_in , 
        \local_node[12].data_out , \local_node[13].clk , 
        \local_node[13].buffer_full_in , \local_node[13].buffer_full_out , 
        \local_node[13].receiving_data , \local_node[13].sending_data , 
        \local_node[13].data_in , \local_node[13].data_out , 
        \local_node[14].clk , \local_node[14].buffer_full_in , 
        \local_node[14].buffer_full_out , \local_node[14].receiving_data , 
        \local_node[14].sending_data , \local_node[14].data_in , 
        \local_node[14].data_out , \local_node[15].clk , 
        \local_node[15].buffer_full_in , \local_node[15].buffer_full_out , 
        \local_node[15].receiving_data , \local_node[15].sending_data , 
        \local_node[15].data_in , \local_node[15].data_out  );
  inout [15:0] \local_node[0].data_in ;
  inout [15:0] \local_node[0].data_out ;
  inout [15:0] \local_node[1].data_in ;
  inout [15:0] \local_node[1].data_out ;
  inout [15:0] \local_node[2].data_in ;
  inout [15:0] \local_node[2].data_out ;
  inout [15:0] \local_node[3].data_in ;
  inout [15:0] \local_node[3].data_out ;
  inout [15:0] \local_node[4].data_in ;
  inout [15:0] \local_node[4].data_out ;
  inout [15:0] \local_node[5].data_in ;
  inout [15:0] \local_node[5].data_out ;
  inout [15:0] \local_node[6].data_in ;
  inout [15:0] \local_node[6].data_out ;
  inout [15:0] \local_node[7].data_in ;
  inout [15:0] \local_node[7].data_out ;
  inout [15:0] \local_node[8].data_in ;
  inout [15:0] \local_node[8].data_out ;
  inout [15:0] \local_node[9].data_in ;
  inout [15:0] \local_node[9].data_out ;
  inout [15:0] \local_node[10].data_in ;
  inout [15:0] \local_node[10].data_out ;
  inout [15:0] \local_node[11].data_in ;
  inout [15:0] \local_node[11].data_out ;
  inout [15:0] \local_node[12].data_in ;
  inout [15:0] \local_node[12].data_out ;
  inout [15:0] \local_node[13].data_in ;
  inout [15:0] \local_node[13].data_out ;
  inout [15:0] \local_node[14].data_in ;
  inout [15:0] \local_node[14].data_out ;
  inout [15:0] \local_node[15].data_in ;
  inout [15:0] \local_node[15].data_out ;
  input \clk.clk , \reset.reset , \local_node[0].clk , \local_node[1].clk ,
         \local_node[2].clk , \local_node[3].clk , \local_node[4].clk ,
         \local_node[5].clk , \local_node[6].clk , \local_node[7].clk ,
         \local_node[8].clk , \local_node[9].clk , \local_node[10].clk ,
         \local_node[11].clk , \local_node[12].clk , \local_node[13].clk ,
         \local_node[14].clk , \local_node[15].clk ;
  inout \local_node[0].buffer_full_in ,  \local_node[0].buffer_full_out , 
     \local_node[0].receiving_data ,  \local_node[0].sending_data , 
     \local_node[1].buffer_full_in ,  \local_node[1].buffer_full_out , 
     \local_node[1].receiving_data ,  \local_node[1].sending_data , 
     \local_node[2].buffer_full_in ,  \local_node[2].buffer_full_out , 
     \local_node[2].receiving_data ,  \local_node[2].sending_data , 
     \local_node[3].buffer_full_in ,  \local_node[3].buffer_full_out , 
     \local_node[3].receiving_data ,  \local_node[3].sending_data , 
     \local_node[4].buffer_full_in ,  \local_node[4].buffer_full_out , 
     \local_node[4].receiving_data ,  \local_node[4].sending_data , 
     \local_node[5].buffer_full_in ,  \local_node[5].buffer_full_out , 
     \local_node[5].receiving_data ,  \local_node[5].sending_data , 
     \local_node[6].buffer_full_in ,  \local_node[6].buffer_full_out , 
     \local_node[6].receiving_data ,  \local_node[6].sending_data , 
     \local_node[7].buffer_full_in ,  \local_node[7].buffer_full_out , 
     \local_node[7].receiving_data ,  \local_node[7].sending_data , 
     \local_node[8].buffer_full_in ,  \local_node[8].buffer_full_out , 
     \local_node[8].receiving_data ,  \local_node[8].sending_data , 
     \local_node[9].buffer_full_in ,  \local_node[9].buffer_full_out , 
     \local_node[9].receiving_data ,  \local_node[9].sending_data , 
     \local_node[10].buffer_full_in ,  \local_node[10].buffer_full_out , 
     \local_node[10].receiving_data ,  \local_node[10].sending_data , 
     \local_node[11].buffer_full_in ,  \local_node[11].buffer_full_out , 
     \local_node[11].receiving_data ,  \local_node[11].sending_data , 
     \local_node[12].buffer_full_in ,  \local_node[12].buffer_full_out , 
     \local_node[12].receiving_data ,  \local_node[12].sending_data , 
     \local_node[13].buffer_full_in ,  \local_node[13].buffer_full_out , 
     \local_node[13].receiving_data ,  \local_node[13].sending_data , 
     \local_node[14].buffer_full_in ,  \local_node[14].buffer_full_out , 
     \local_node[14].receiving_data ,  \local_node[14].sending_data , 
     \local_node[15].buffer_full_in ,  \local_node[15].buffer_full_out , 
     \local_node[15].receiving_data ,  \local_node[15].sending_data ;
  wire   \local_node[16].clk ;
  tri   \local_node[0].buffer_full_in ;
  tri   \local_node[0].buffer_full_out ;
  tri   \local_node[0].receiving_data ;
  tri   \local_node[0].sending_data ;
  tri   \local_node[0].data_in[15] ;
  tri   \local_node[0].data_in[14] ;
  tri   \local_node[0].data_in[13] ;
  tri   \local_node[0].data_in[12] ;
  tri   \local_node[0].data_in[11] ;
  tri   \local_node[0].data_in[10] ;
  tri   \local_node[0].data_in[9] ;
  tri   \local_node[0].data_in[8] ;
  tri   \local_node[0].data_in[7] ;
  tri   \local_node[0].data_in[6] ;
  tri   \local_node[0].data_in[5] ;
  tri   \local_node[0].data_in[4] ;
  tri   \local_node[0].data_in[3] ;
  tri   \local_node[0].data_in[2] ;
  tri   \local_node[0].data_in[1] ;
  tri   \local_node[0].data_in[0] ;
  tri   \local_node[0].data_out[15] ;
  tri   \local_node[0].data_out[14] ;
  tri   \local_node[0].data_out[13] ;
  tri   \local_node[0].data_out[12] ;
  tri   \local_node[0].data_out[11] ;
  tri   \local_node[0].data_out[10] ;
  tri   \local_node[0].data_out[9] ;
  tri   \local_node[0].data_out[8] ;
  tri   \local_node[0].data_out[7] ;
  tri   \local_node[0].data_out[6] ;
  tri   \local_node[0].data_out[5] ;
  tri   \local_node[0].data_out[4] ;
  tri   \local_node[0].data_out[3] ;
  tri   \local_node[0].data_out[2] ;
  tri   \local_node[0].data_out[1] ;
  tri   \local_node[0].data_out[0] ;
  tri   \local_node[1].buffer_full_in ;
  tri   \local_node[1].buffer_full_out ;
  tri   \local_node[1].receiving_data ;
  tri   \local_node[1].sending_data ;
  tri   \local_node[1].data_in[15] ;
  tri   \local_node[1].data_in[14] ;
  tri   \local_node[1].data_in[13] ;
  tri   \local_node[1].data_in[12] ;
  tri   \local_node[1].data_in[11] ;
  tri   \local_node[1].data_in[10] ;
  tri   \local_node[1].data_in[9] ;
  tri   \local_node[1].data_in[8] ;
  tri   \local_node[1].data_in[7] ;
  tri   \local_node[1].data_in[6] ;
  tri   \local_node[1].data_in[5] ;
  tri   \local_node[1].data_in[4] ;
  tri   \local_node[1].data_in[3] ;
  tri   \local_node[1].data_in[2] ;
  tri   \local_node[1].data_in[1] ;
  tri   \local_node[1].data_in[0] ;
  tri   \local_node[1].data_out[15] ;
  tri   \local_node[1].data_out[14] ;
  tri   \local_node[1].data_out[13] ;
  tri   \local_node[1].data_out[12] ;
  tri   \local_node[1].data_out[11] ;
  tri   \local_node[1].data_out[10] ;
  tri   \local_node[1].data_out[9] ;
  tri   \local_node[1].data_out[8] ;
  tri   \local_node[1].data_out[7] ;
  tri   \local_node[1].data_out[6] ;
  tri   \local_node[1].data_out[5] ;
  tri   \local_node[1].data_out[4] ;
  tri   \local_node[1].data_out[3] ;
  tri   \local_node[1].data_out[2] ;
  tri   \local_node[1].data_out[1] ;
  tri   \local_node[1].data_out[0] ;
  tri   \local_node[2].buffer_full_in ;
  tri   \local_node[2].buffer_full_out ;
  tri   \local_node[2].receiving_data ;
  tri   \local_node[2].sending_data ;
  tri   \local_node[2].data_in[15] ;
  tri   \local_node[2].data_in[14] ;
  tri   \local_node[2].data_in[13] ;
  tri   \local_node[2].data_in[12] ;
  tri   \local_node[2].data_in[11] ;
  tri   \local_node[2].data_in[10] ;
  tri   \local_node[2].data_in[9] ;
  tri   \local_node[2].data_in[8] ;
  tri   \local_node[2].data_in[7] ;
  tri   \local_node[2].data_in[6] ;
  tri   \local_node[2].data_in[5] ;
  tri   \local_node[2].data_in[4] ;
  tri   \local_node[2].data_in[3] ;
  tri   \local_node[2].data_in[2] ;
  tri   \local_node[2].data_in[1] ;
  tri   \local_node[2].data_in[0] ;
  tri   \local_node[2].data_out[15] ;
  tri   \local_node[2].data_out[14] ;
  tri   \local_node[2].data_out[13] ;
  tri   \local_node[2].data_out[12] ;
  tri   \local_node[2].data_out[11] ;
  tri   \local_node[2].data_out[10] ;
  tri   \local_node[2].data_out[9] ;
  tri   \local_node[2].data_out[8] ;
  tri   \local_node[2].data_out[7] ;
  tri   \local_node[2].data_out[6] ;
  tri   \local_node[2].data_out[5] ;
  tri   \local_node[2].data_out[4] ;
  tri   \local_node[2].data_out[3] ;
  tri   \local_node[2].data_out[2] ;
  tri   \local_node[2].data_out[1] ;
  tri   \local_node[2].data_out[0] ;
  tri   \local_node[3].buffer_full_in ;
  tri   \local_node[3].buffer_full_out ;
  tri   \local_node[3].receiving_data ;
  tri   \local_node[3].sending_data ;
  tri   \local_node[3].data_in[15] ;
  tri   \local_node[3].data_in[14] ;
  tri   \local_node[3].data_in[13] ;
  tri   \local_node[3].data_in[12] ;
  tri   \local_node[3].data_in[11] ;
  tri   \local_node[3].data_in[10] ;
  tri   \local_node[3].data_in[9] ;
  tri   \local_node[3].data_in[8] ;
  tri   \local_node[3].data_in[7] ;
  tri   \local_node[3].data_in[6] ;
  tri   \local_node[3].data_in[5] ;
  tri   \local_node[3].data_in[4] ;
  tri   \local_node[3].data_in[3] ;
  tri   \local_node[3].data_in[2] ;
  tri   \local_node[3].data_in[1] ;
  tri   \local_node[3].data_in[0] ;
  tri   \local_node[3].data_out[15] ;
  tri   \local_node[3].data_out[14] ;
  tri   \local_node[3].data_out[13] ;
  tri   \local_node[3].data_out[12] ;
  tri   \local_node[3].data_out[11] ;
  tri   \local_node[3].data_out[10] ;
  tri   \local_node[3].data_out[9] ;
  tri   \local_node[3].data_out[8] ;
  tri   \local_node[3].data_out[7] ;
  tri   \local_node[3].data_out[6] ;
  tri   \local_node[3].data_out[5] ;
  tri   \local_node[3].data_out[4] ;
  tri   \local_node[3].data_out[3] ;
  tri   \local_node[3].data_out[2] ;
  tri   \local_node[3].data_out[1] ;
  tri   \local_node[3].data_out[0] ;
  tri   \local_node[4].buffer_full_in ;
  tri   \local_node[4].buffer_full_out ;
  tri   \local_node[4].receiving_data ;
  tri   \local_node[4].sending_data ;
  tri   \local_node[4].data_in[15] ;
  tri   \local_node[4].data_in[14] ;
  tri   \local_node[4].data_in[13] ;
  tri   \local_node[4].data_in[12] ;
  tri   \local_node[4].data_in[11] ;
  tri   \local_node[4].data_in[10] ;
  tri   \local_node[4].data_in[9] ;
  tri   \local_node[4].data_in[8] ;
  tri   \local_node[4].data_in[7] ;
  tri   \local_node[4].data_in[6] ;
  tri   \local_node[4].data_in[5] ;
  tri   \local_node[4].data_in[4] ;
  tri   \local_node[4].data_in[3] ;
  tri   \local_node[4].data_in[2] ;
  tri   \local_node[4].data_in[1] ;
  tri   \local_node[4].data_in[0] ;
  tri   \local_node[4].data_out[15] ;
  tri   \local_node[4].data_out[14] ;
  tri   \local_node[4].data_out[13] ;
  tri   \local_node[4].data_out[12] ;
  tri   \local_node[4].data_out[11] ;
  tri   \local_node[4].data_out[10] ;
  tri   \local_node[4].data_out[9] ;
  tri   \local_node[4].data_out[8] ;
  tri   \local_node[4].data_out[7] ;
  tri   \local_node[4].data_out[6] ;
  tri   \local_node[4].data_out[5] ;
  tri   \local_node[4].data_out[4] ;
  tri   \local_node[4].data_out[3] ;
  tri   \local_node[4].data_out[2] ;
  tri   \local_node[4].data_out[1] ;
  tri   \local_node[4].data_out[0] ;
  tri   \local_node[5].buffer_full_in ;
  tri   \local_node[5].buffer_full_out ;
  tri   \local_node[5].receiving_data ;
  tri   \local_node[5].sending_data ;
  tri   \local_node[5].data_in[15] ;
  tri   \local_node[5].data_in[14] ;
  tri   \local_node[5].data_in[13] ;
  tri   \local_node[5].data_in[12] ;
  tri   \local_node[5].data_in[11] ;
  tri   \local_node[5].data_in[10] ;
  tri   \local_node[5].data_in[9] ;
  tri   \local_node[5].data_in[8] ;
  tri   \local_node[5].data_in[7] ;
  tri   \local_node[5].data_in[6] ;
  tri   \local_node[5].data_in[5] ;
  tri   \local_node[5].data_in[4] ;
  tri   \local_node[5].data_in[3] ;
  tri   \local_node[5].data_in[2] ;
  tri   \local_node[5].data_in[1] ;
  tri   \local_node[5].data_in[0] ;
  tri   \local_node[5].data_out[15] ;
  tri   \local_node[5].data_out[14] ;
  tri   \local_node[5].data_out[13] ;
  tri   \local_node[5].data_out[12] ;
  tri   \local_node[5].data_out[11] ;
  tri   \local_node[5].data_out[10] ;
  tri   \local_node[5].data_out[9] ;
  tri   \local_node[5].data_out[8] ;
  tri   \local_node[5].data_out[7] ;
  tri   \local_node[5].data_out[6] ;
  tri   \local_node[5].data_out[5] ;
  tri   \local_node[5].data_out[4] ;
  tri   \local_node[5].data_out[3] ;
  tri   \local_node[5].data_out[2] ;
  tri   \local_node[5].data_out[1] ;
  tri   \local_node[5].data_out[0] ;
  tri   \local_node[6].buffer_full_in ;
  tri   \local_node[6].buffer_full_out ;
  tri   \local_node[6].receiving_data ;
  tri   \local_node[6].sending_data ;
  tri   \local_node[6].data_in[15] ;
  tri   \local_node[6].data_in[14] ;
  tri   \local_node[6].data_in[13] ;
  tri   \local_node[6].data_in[12] ;
  tri   \local_node[6].data_in[11] ;
  tri   \local_node[6].data_in[10] ;
  tri   \local_node[6].data_in[9] ;
  tri   \local_node[6].data_in[8] ;
  tri   \local_node[6].data_in[7] ;
  tri   \local_node[6].data_in[6] ;
  tri   \local_node[6].data_in[5] ;
  tri   \local_node[6].data_in[4] ;
  tri   \local_node[6].data_in[3] ;
  tri   \local_node[6].data_in[2] ;
  tri   \local_node[6].data_in[1] ;
  tri   \local_node[6].data_in[0] ;
  tri   \local_node[6].data_out[15] ;
  tri   \local_node[6].data_out[14] ;
  tri   \local_node[6].data_out[13] ;
  tri   \local_node[6].data_out[12] ;
  tri   \local_node[6].data_out[11] ;
  tri   \local_node[6].data_out[10] ;
  tri   \local_node[6].data_out[9] ;
  tri   \local_node[6].data_out[8] ;
  tri   \local_node[6].data_out[7] ;
  tri   \local_node[6].data_out[6] ;
  tri   \local_node[6].data_out[5] ;
  tri   \local_node[6].data_out[4] ;
  tri   \local_node[6].data_out[3] ;
  tri   \local_node[6].data_out[2] ;
  tri   \local_node[6].data_out[1] ;
  tri   \local_node[6].data_out[0] ;
  tri   \local_node[7].buffer_full_in ;
  tri   \local_node[7].buffer_full_out ;
  tri   \local_node[7].receiving_data ;
  tri   \local_node[7].sending_data ;
  tri   \local_node[7].data_in[15] ;
  tri   \local_node[7].data_in[14] ;
  tri   \local_node[7].data_in[13] ;
  tri   \local_node[7].data_in[12] ;
  tri   \local_node[7].data_in[11] ;
  tri   \local_node[7].data_in[10] ;
  tri   \local_node[7].data_in[9] ;
  tri   \local_node[7].data_in[8] ;
  tri   \local_node[7].data_in[7] ;
  tri   \local_node[7].data_in[6] ;
  tri   \local_node[7].data_in[5] ;
  tri   \local_node[7].data_in[4] ;
  tri   \local_node[7].data_in[3] ;
  tri   \local_node[7].data_in[2] ;
  tri   \local_node[7].data_in[1] ;
  tri   \local_node[7].data_in[0] ;
  tri   \local_node[7].data_out[15] ;
  tri   \local_node[7].data_out[14] ;
  tri   \local_node[7].data_out[13] ;
  tri   \local_node[7].data_out[12] ;
  tri   \local_node[7].data_out[11] ;
  tri   \local_node[7].data_out[10] ;
  tri   \local_node[7].data_out[9] ;
  tri   \local_node[7].data_out[8] ;
  tri   \local_node[7].data_out[7] ;
  tri   \local_node[7].data_out[6] ;
  tri   \local_node[7].data_out[5] ;
  tri   \local_node[7].data_out[4] ;
  tri   \local_node[7].data_out[3] ;
  tri   \local_node[7].data_out[2] ;
  tri   \local_node[7].data_out[1] ;
  tri   \local_node[7].data_out[0] ;
  tri   \local_node[8].buffer_full_in ;
  tri   \local_node[8].buffer_full_out ;
  tri   \local_node[8].receiving_data ;
  tri   \local_node[8].sending_data ;
  tri   \local_node[8].data_in[15] ;
  tri   \local_node[8].data_in[14] ;
  tri   \local_node[8].data_in[13] ;
  tri   \local_node[8].data_in[12] ;
  tri   \local_node[8].data_in[11] ;
  tri   \local_node[8].data_in[10] ;
  tri   \local_node[8].data_in[9] ;
  tri   \local_node[8].data_in[8] ;
  tri   \local_node[8].data_in[7] ;
  tri   \local_node[8].data_in[6] ;
  tri   \local_node[8].data_in[5] ;
  tri   \local_node[8].data_in[4] ;
  tri   \local_node[8].data_in[3] ;
  tri   \local_node[8].data_in[2] ;
  tri   \local_node[8].data_in[1] ;
  tri   \local_node[8].data_in[0] ;
  tri   \local_node[8].data_out[15] ;
  tri   \local_node[8].data_out[14] ;
  tri   \local_node[8].data_out[13] ;
  tri   \local_node[8].data_out[12] ;
  tri   \local_node[8].data_out[11] ;
  tri   \local_node[8].data_out[10] ;
  tri   \local_node[8].data_out[9] ;
  tri   \local_node[8].data_out[8] ;
  tri   \local_node[8].data_out[7] ;
  tri   \local_node[8].data_out[6] ;
  tri   \local_node[8].data_out[5] ;
  tri   \local_node[8].data_out[4] ;
  tri   \local_node[8].data_out[3] ;
  tri   \local_node[8].data_out[2] ;
  tri   \local_node[8].data_out[1] ;
  tri   \local_node[8].data_out[0] ;
  tri   \local_node[9].buffer_full_in ;
  tri   \local_node[9].buffer_full_out ;
  tri   \local_node[9].receiving_data ;
  tri   \local_node[9].sending_data ;
  tri   \local_node[9].data_in[15] ;
  tri   \local_node[9].data_in[14] ;
  tri   \local_node[9].data_in[13] ;
  tri   \local_node[9].data_in[12] ;
  tri   \local_node[9].data_in[11] ;
  tri   \local_node[9].data_in[10] ;
  tri   \local_node[9].data_in[9] ;
  tri   \local_node[9].data_in[8] ;
  tri   \local_node[9].data_in[7] ;
  tri   \local_node[9].data_in[6] ;
  tri   \local_node[9].data_in[5] ;
  tri   \local_node[9].data_in[4] ;
  tri   \local_node[9].data_in[3] ;
  tri   \local_node[9].data_in[2] ;
  tri   \local_node[9].data_in[1] ;
  tri   \local_node[9].data_in[0] ;
  tri   \local_node[9].data_out[15] ;
  tri   \local_node[9].data_out[14] ;
  tri   \local_node[9].data_out[13] ;
  tri   \local_node[9].data_out[12] ;
  tri   \local_node[9].data_out[11] ;
  tri   \local_node[9].data_out[10] ;
  tri   \local_node[9].data_out[9] ;
  tri   \local_node[9].data_out[8] ;
  tri   \local_node[9].data_out[7] ;
  tri   \local_node[9].data_out[6] ;
  tri   \local_node[9].data_out[5] ;
  tri   \local_node[9].data_out[4] ;
  tri   \local_node[9].data_out[3] ;
  tri   \local_node[9].data_out[2] ;
  tri   \local_node[9].data_out[1] ;
  tri   \local_node[9].data_out[0] ;
  tri   \local_node[10].buffer_full_in ;
  tri   \local_node[10].buffer_full_out ;
  tri   \local_node[10].receiving_data ;
  tri   \local_node[10].sending_data ;
  tri   \local_node[10].data_in[15] ;
  tri   \local_node[10].data_in[14] ;
  tri   \local_node[10].data_in[13] ;
  tri   \local_node[10].data_in[12] ;
  tri   \local_node[10].data_in[11] ;
  tri   \local_node[10].data_in[10] ;
  tri   \local_node[10].data_in[9] ;
  tri   \local_node[10].data_in[8] ;
  tri   \local_node[10].data_in[7] ;
  tri   \local_node[10].data_in[6] ;
  tri   \local_node[10].data_in[5] ;
  tri   \local_node[10].data_in[4] ;
  tri   \local_node[10].data_in[3] ;
  tri   \local_node[10].data_in[2] ;
  tri   \local_node[10].data_in[1] ;
  tri   \local_node[10].data_in[0] ;
  tri   \local_node[10].data_out[15] ;
  tri   \local_node[10].data_out[14] ;
  tri   \local_node[10].data_out[13] ;
  tri   \local_node[10].data_out[12] ;
  tri   \local_node[10].data_out[11] ;
  tri   \local_node[10].data_out[10] ;
  tri   \local_node[10].data_out[9] ;
  tri   \local_node[10].data_out[8] ;
  tri   \local_node[10].data_out[7] ;
  tri   \local_node[10].data_out[6] ;
  tri   \local_node[10].data_out[5] ;
  tri   \local_node[10].data_out[4] ;
  tri   \local_node[10].data_out[3] ;
  tri   \local_node[10].data_out[2] ;
  tri   \local_node[10].data_out[1] ;
  tri   \local_node[10].data_out[0] ;
  tri   \local_node[11].buffer_full_in ;
  tri   \local_node[11].buffer_full_out ;
  tri   \local_node[11].receiving_data ;
  tri   \local_node[11].sending_data ;
  tri   \local_node[11].data_in[15] ;
  tri   \local_node[11].data_in[14] ;
  tri   \local_node[11].data_in[13] ;
  tri   \local_node[11].data_in[12] ;
  tri   \local_node[11].data_in[11] ;
  tri   \local_node[11].data_in[10] ;
  tri   \local_node[11].data_in[9] ;
  tri   \local_node[11].data_in[8] ;
  tri   \local_node[11].data_in[7] ;
  tri   \local_node[11].data_in[6] ;
  tri   \local_node[11].data_in[5] ;
  tri   \local_node[11].data_in[4] ;
  tri   \local_node[11].data_in[3] ;
  tri   \local_node[11].data_in[2] ;
  tri   \local_node[11].data_in[1] ;
  tri   \local_node[11].data_in[0] ;
  tri   \local_node[11].data_out[15] ;
  tri   \local_node[11].data_out[14] ;
  tri   \local_node[11].data_out[13] ;
  tri   \local_node[11].data_out[12] ;
  tri   \local_node[11].data_out[11] ;
  tri   \local_node[11].data_out[10] ;
  tri   \local_node[11].data_out[9] ;
  tri   \local_node[11].data_out[8] ;
  tri   \local_node[11].data_out[7] ;
  tri   \local_node[11].data_out[6] ;
  tri   \local_node[11].data_out[5] ;
  tri   \local_node[11].data_out[4] ;
  tri   \local_node[11].data_out[3] ;
  tri   \local_node[11].data_out[2] ;
  tri   \local_node[11].data_out[1] ;
  tri   \local_node[11].data_out[0] ;
  tri   \local_node[12].buffer_full_in ;
  tri   \local_node[12].buffer_full_out ;
  tri   \local_node[12].receiving_data ;
  tri   \local_node[12].sending_data ;
  tri   \local_node[12].data_in[15] ;
  tri   \local_node[12].data_in[14] ;
  tri   \local_node[12].data_in[13] ;
  tri   \local_node[12].data_in[12] ;
  tri   \local_node[12].data_in[11] ;
  tri   \local_node[12].data_in[10] ;
  tri   \local_node[12].data_in[9] ;
  tri   \local_node[12].data_in[8] ;
  tri   \local_node[12].data_in[7] ;
  tri   \local_node[12].data_in[6] ;
  tri   \local_node[12].data_in[5] ;
  tri   \local_node[12].data_in[4] ;
  tri   \local_node[12].data_in[3] ;
  tri   \local_node[12].data_in[2] ;
  tri   \local_node[12].data_in[1] ;
  tri   \local_node[12].data_in[0] ;
  tri   \local_node[12].data_out[15] ;
  tri   \local_node[12].data_out[14] ;
  tri   \local_node[12].data_out[13] ;
  tri   \local_node[12].data_out[12] ;
  tri   \local_node[12].data_out[11] ;
  tri   \local_node[12].data_out[10] ;
  tri   \local_node[12].data_out[9] ;
  tri   \local_node[12].data_out[8] ;
  tri   \local_node[12].data_out[7] ;
  tri   \local_node[12].data_out[6] ;
  tri   \local_node[12].data_out[5] ;
  tri   \local_node[12].data_out[4] ;
  tri   \local_node[12].data_out[3] ;
  tri   \local_node[12].data_out[2] ;
  tri   \local_node[12].data_out[1] ;
  tri   \local_node[12].data_out[0] ;
  tri   \local_node[13].buffer_full_in ;
  tri   \local_node[13].buffer_full_out ;
  tri   \local_node[13].receiving_data ;
  tri   \local_node[13].sending_data ;
  tri   \local_node[13].data_in[15] ;
  tri   \local_node[13].data_in[14] ;
  tri   \local_node[13].data_in[13] ;
  tri   \local_node[13].data_in[12] ;
  tri   \local_node[13].data_in[11] ;
  tri   \local_node[13].data_in[10] ;
  tri   \local_node[13].data_in[9] ;
  tri   \local_node[13].data_in[8] ;
  tri   \local_node[13].data_in[7] ;
  tri   \local_node[13].data_in[6] ;
  tri   \local_node[13].data_in[5] ;
  tri   \local_node[13].data_in[4] ;
  tri   \local_node[13].data_in[3] ;
  tri   \local_node[13].data_in[2] ;
  tri   \local_node[13].data_in[1] ;
  tri   \local_node[13].data_in[0] ;
  tri   \local_node[13].data_out[15] ;
  tri   \local_node[13].data_out[14] ;
  tri   \local_node[13].data_out[13] ;
  tri   \local_node[13].data_out[12] ;
  tri   \local_node[13].data_out[11] ;
  tri   \local_node[13].data_out[10] ;
  tri   \local_node[13].data_out[9] ;
  tri   \local_node[13].data_out[8] ;
  tri   \local_node[13].data_out[7] ;
  tri   \local_node[13].data_out[6] ;
  tri   \local_node[13].data_out[5] ;
  tri   \local_node[13].data_out[4] ;
  tri   \local_node[13].data_out[3] ;
  tri   \local_node[13].data_out[2] ;
  tri   \local_node[13].data_out[1] ;
  tri   \local_node[13].data_out[0] ;
  tri   \local_node[14].buffer_full_in ;
  tri   \local_node[14].buffer_full_out ;
  tri   \local_node[14].receiving_data ;
  tri   \local_node[14].sending_data ;
  tri   \local_node[14].data_in[15] ;
  tri   \local_node[14].data_in[14] ;
  tri   \local_node[14].data_in[13] ;
  tri   \local_node[14].data_in[12] ;
  tri   \local_node[14].data_in[11] ;
  tri   \local_node[14].data_in[10] ;
  tri   \local_node[14].data_in[9] ;
  tri   \local_node[14].data_in[8] ;
  tri   \local_node[14].data_in[7] ;
  tri   \local_node[14].data_in[6] ;
  tri   \local_node[14].data_in[5] ;
  tri   \local_node[14].data_in[4] ;
  tri   \local_node[14].data_in[3] ;
  tri   \local_node[14].data_in[2] ;
  tri   \local_node[14].data_in[1] ;
  tri   \local_node[14].data_in[0] ;
  tri   \local_node[14].data_out[15] ;
  tri   \local_node[14].data_out[14] ;
  tri   \local_node[14].data_out[13] ;
  tri   \local_node[14].data_out[12] ;
  tri   \local_node[14].data_out[11] ;
  tri   \local_node[14].data_out[10] ;
  tri   \local_node[14].data_out[9] ;
  tri   \local_node[14].data_out[8] ;
  tri   \local_node[14].data_out[7] ;
  tri   \local_node[14].data_out[6] ;
  tri   \local_node[14].data_out[5] ;
  tri   \local_node[14].data_out[4] ;
  tri   \local_node[14].data_out[3] ;
  tri   \local_node[14].data_out[2] ;
  tri   \local_node[14].data_out[1] ;
  tri   \local_node[14].data_out[0] ;
  tri   \local_node[16].buffer_full_in ;
  tri   \local_node[16].buffer_full_out ;
  tri   \local_node[16].receiving_data ;
  tri   \local_node[16].sending_data ;
  tri   \local_node[16].data_in[15] ;
  tri   \local_node[16].data_in[14] ;
  tri   \local_node[16].data_in[13] ;
  tri   \local_node[16].data_in[12] ;
  tri   \local_node[16].data_in[11] ;
  tri   \local_node[16].data_in[10] ;
  tri   \local_node[16].data_in[9] ;
  tri   \local_node[16].data_in[8] ;
  tri   \local_node[16].data_in[7] ;
  tri   \local_node[16].data_in[6] ;
  tri   \local_node[16].data_in[5] ;
  tri   \local_node[16].data_in[4] ;
  tri   \local_node[16].data_in[3] ;
  tri   \local_node[16].data_in[2] ;
  tri   \local_node[16].data_in[1] ;
  tri   \local_node[16].data_in[0] ;
  tri   \local_node[16].data_out[15] ;
  tri   \local_node[16].data_out[14] ;
  tri   \local_node[16].data_out[13] ;
  tri   \local_node[16].data_out[12] ;
  tri   \local_node[16].data_out[11] ;
  tri   \local_node[16].data_out[10] ;
  tri   \local_node[16].data_out[9] ;
  tri   \local_node[16].data_out[8] ;
  tri   \local_node[16].data_out[7] ;
  tri   \local_node[16].data_out[6] ;
  tri   \local_node[16].data_out[5] ;
  tri   \local_node[16].data_out[4] ;
  tri   \local_node[16].data_out[3] ;
  tri   \local_node[16].data_out[2] ;
  tri   \local_node[16].data_out[1] ;
  tri   \local_node[16].data_out[0] ;
  assign \local_node[16].clk  = \local_node[15].clk ;
  tran( \local_node[16].buffer_full_in , \local_node[15].buffer_full_in );
  tran( \local_node[16].buffer_full_out , \local_node[15].buffer_full_out );
  tran( \local_node[16].receiving_data , \local_node[15].receiving_data );
  tran( \local_node[16].sending_data , \local_node[15].sending_data );
  tran( \local_node[16].data_in[15] , \local_node[15].data_in  [15]);
  tran( \local_node[16].data_in[14] , \local_node[15].data_in  [14]);
  tran( \local_node[16].data_in[13] , \local_node[15].data_in  [13]);
  tran( \local_node[16].data_in[12] , \local_node[15].data_in  [12]);
  tran( \local_node[16].data_in[11] , \local_node[15].data_in  [11]);
  tran( \local_node[16].data_in[10] , \local_node[15].data_in  [10]);
  tran( \local_node[16].data_in[9] , \local_node[15].data_in  [9]);
  tran( \local_node[16].data_in[8] , \local_node[15].data_in  [8]);
  tran( \local_node[16].data_in[7] , \local_node[15].data_in  [7]);
  tran( \local_node[16].data_in[6] , \local_node[15].data_in  [6]);
  tran( \local_node[16].data_in[5] , \local_node[15].data_in  [5]);
  tran( \local_node[16].data_in[4] , \local_node[15].data_in  [4]);
  tran( \local_node[16].data_in[3] , \local_node[15].data_in  [3]);
  tran( \local_node[16].data_in[2] , \local_node[15].data_in  [2]);
  tran( \local_node[16].data_in[1] , \local_node[15].data_in  [1]);
  tran( \local_node[16].data_in[0] , \local_node[15].data_in  [0]);
  tran( \local_node[16].data_out[15] , \local_node[15].data_out  [15]);
  tran( \local_node[16].data_out[14] , \local_node[15].data_out  [14]);
  tran( \local_node[16].data_out[13] , \local_node[15].data_out  [13]);
  tran( \local_node[16].data_out[12] , \local_node[15].data_out  [12]);
  tran( \local_node[16].data_out[11] , \local_node[15].data_out  [11]);
  tran( \local_node[16].data_out[10] , \local_node[15].data_out  [10]);
  tran( \local_node[16].data_out[9] , \local_node[15].data_out  [9]);
  tran( \local_node[16].data_out[8] , \local_node[15].data_out  [8]);
  tran( \local_node[16].data_out[7] , \local_node[15].data_out  [7]);
  tran( \local_node[16].data_out[6] , \local_node[15].data_out  [6]);
  tran( \local_node[16].data_out[5] , \local_node[15].data_out  [5]);
  tran( \local_node[16].data_out[4] , \local_node[15].data_out  [4]);
  tran( \local_node[16].data_out[3] , \local_node[15].data_out  [3]);
  tran( \local_node[16].data_out[2] , \local_node[15].data_out  [2]);
  tran( \local_node[16].data_out[1] , \local_node[15].data_out  [1]);
  tran( \local_node[16].data_out[0] , \local_node[15].data_out  [0]);

  node3_NODE_X0_NODE_Y0I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__ tl ( 
        .\clk.clk (\clk.clk ), .\reset.reset (\reset.reset ), 
        .\local_node.clk (\local_node[0].clk ), .\local_node.buffer_full_in (
        \local_node[0].buffer_full_in ), .\local_node.buffer_full_out (
        \local_node[0].buffer_full_out ), .\local_node.receiving_data (
        \local_node[0].receiving_data ), .\local_node.sending_data (
        \local_node[0].sending_data ), .\local_node.data_in ({
        \local_node[0].data_in  [15], \local_node[0].data_in  [14], 
        \local_node[0].data_in  [13], \local_node[0].data_in  [12], 
        \local_node[0].data_in  [11], \local_node[0].data_in  [10], 
        \local_node[0].data_in  [9], \local_node[0].data_in  [8], 
        \local_node[0].data_in  [7], \local_node[0].data_in  [6], 
        \local_node[0].data_in  [5], \local_node[0].data_in  [4], 
        \local_node[0].data_in  [3], \local_node[0].data_in  [2], 
        \local_node[0].data_in  [1], \local_node[0].data_in  [0]}), 
        .\local_node.data_out ({\local_node[0].data_out  [15], 
        \local_node[0].data_out  [14], \local_node[0].data_out  [13], 
        \local_node[0].data_out  [12], \local_node[0].data_out  [11], 
        \local_node[0].data_out  [10], \local_node[0].data_out  [9], 
        \local_node[0].data_out  [8], \local_node[0].data_out  [7], 
        \local_node[0].data_out  [6], \local_node[0].data_out  [5], 
        \local_node[0].data_out  [4], \local_node[0].data_out  [3], 
        \local_node[0].data_out  [2], \local_node[0].data_out  [1], 
        \local_node[0].data_out  [0]}), .\node_0.clk (\clk.clk ), 
        .\node_0.buffer_full_in (1'b0), .\node_0.receiving_data (1'b0), 
        .\node_0.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_1.clk (
        \clk.clk ), .\node_1.buffer_full_in (1'b0), .\node_1.receiving_data (
        1'b0), .\node_1.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  node3_NODE_X3_NODE_Y0I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__ tr ( 
        .\clk.clk (\clk.clk ), .\reset.reset (\reset.reset ), 
        .\local_node.clk (\local_node[3].clk ), .\local_node.buffer_full_in (
        \local_node[3].buffer_full_in ), .\local_node.buffer_full_out (
        \local_node[3].buffer_full_out ), .\local_node.receiving_data (
        \local_node[3].receiving_data ), .\local_node.sending_data (
        \local_node[3].sending_data ), .\local_node.data_in ({
        \local_node[3].data_in  [15], \local_node[3].data_in  [14], 
        \local_node[3].data_in  [13], \local_node[3].data_in  [12], 
        \local_node[3].data_in  [11], \local_node[3].data_in  [10], 
        \local_node[3].data_in  [9], \local_node[3].data_in  [8], 
        \local_node[3].data_in  [7], \local_node[3].data_in  [6], 
        \local_node[3].data_in  [5], \local_node[3].data_in  [4], 
        \local_node[3].data_in  [3], \local_node[3].data_in  [2], 
        \local_node[3].data_in  [1], \local_node[3].data_in  [0]}), 
        .\local_node.data_out ({\local_node[3].data_out  [15], 
        \local_node[3].data_out  [14], \local_node[3].data_out  [13], 
        \local_node[3].data_out  [12], \local_node[3].data_out  [11], 
        \local_node[3].data_out  [10], \local_node[3].data_out  [9], 
        \local_node[3].data_out  [8], \local_node[3].data_out  [7], 
        \local_node[3].data_out  [6], \local_node[3].data_out  [5], 
        \local_node[3].data_out  [4], \local_node[3].data_out  [3], 
        \local_node[3].data_out  [2], \local_node[3].data_out  [1], 
        \local_node[3].data_out  [0]}), .\node_0.clk (\clk.clk ), 
        .\node_0.buffer_full_in (1'b0), .\node_0.receiving_data (1'b0), 
        .\node_0.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_1.clk (
        \clk.clk ), .\node_1.buffer_full_in (1'b0), .\node_1.receiving_data (
        1'b0), .\node_1.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  node3_NODE_X0_NODE_Y3I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__ bl ( 
        .\clk.clk (\clk.clk ), .\reset.reset (\reset.reset ), 
        .\local_node.clk (\local_node[12].clk ), .\local_node.buffer_full_in (
        \local_node[12].buffer_full_in ), .\local_node.buffer_full_out (
        \local_node[12].buffer_full_out ), .\local_node.receiving_data (
        \local_node[12].receiving_data ), .\local_node.sending_data (
        \local_node[12].sending_data ), .\local_node.data_in ({
        \local_node[12].data_in  [15], \local_node[12].data_in  [14], 
        \local_node[12].data_in  [13], \local_node[12].data_in  [12], 
        \local_node[12].data_in  [11], \local_node[12].data_in  [10], 
        \local_node[12].data_in  [9], \local_node[12].data_in  [8], 
        \local_node[12].data_in  [7], \local_node[12].data_in  [6], 
        \local_node[12].data_in  [5], \local_node[12].data_in  [4], 
        \local_node[12].data_in  [3], \local_node[12].data_in  [2], 
        \local_node[12].data_in  [1], \local_node[12].data_in  [0]}), 
        .\local_node.data_out ({\local_node[12].data_out  [15], 
        \local_node[12].data_out  [14], \local_node[12].data_out  [13], 
        \local_node[12].data_out  [12], \local_node[12].data_out  [11], 
        \local_node[12].data_out  [10], \local_node[12].data_out  [9], 
        \local_node[12].data_out  [8], \local_node[12].data_out  [7], 
        \local_node[12].data_out  [6], \local_node[12].data_out  [5], 
        \local_node[12].data_out  [4], \local_node[12].data_out  [3], 
        \local_node[12].data_out  [2], \local_node[12].data_out  [1], 
        \local_node[12].data_out  [0]}), .\node_0.clk (\clk.clk ), 
        .\node_0.buffer_full_in (1'b0), .\node_0.receiving_data (1'b0), 
        .\node_0.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_1.clk (
        \clk.clk ), .\node_1.buffer_full_in (1'b0), .\node_1.receiving_data (
        1'b0), .\node_1.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  node3_NODE_X3_NODE_Y3I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__ br ( 
        .\clk.clk (\clk.clk ), .\reset.reset (\reset.reset ), 
        .\local_node.clk (\local_node[16].clk ), .\local_node.buffer_full_in (
        \local_node[16].buffer_full_in ), .\local_node.buffer_full_out (
        \local_node[16].buffer_full_out ), .\local_node.receiving_data (
        \local_node[16].receiving_data ), .\local_node.sending_data (
        \local_node[16].sending_data ), .\local_node.data_in ({
        \local_node[16].data_in[15] , \local_node[16].data_in[14] , 
        \local_node[16].data_in[13] , \local_node[16].data_in[12] , 
        \local_node[16].data_in[11] , \local_node[16].data_in[10] , 
        \local_node[16].data_in[9] , \local_node[16].data_in[8] , 
        \local_node[16].data_in[7] , \local_node[16].data_in[6] , 
        \local_node[16].data_in[5] , \local_node[16].data_in[4] , 
        \local_node[16].data_in[3] , \local_node[16].data_in[2] , 
        \local_node[16].data_in[1] , \local_node[16].data_in[0] }), 
        .\local_node.data_out ({\local_node[16].data_out[15] , 
        \local_node[16].data_out[14] , \local_node[16].data_out[13] , 
        \local_node[16].data_out[12] , \local_node[16].data_out[11] , 
        \local_node[16].data_out[10] , \local_node[16].data_out[9] , 
        \local_node[16].data_out[8] , \local_node[16].data_out[7] , 
        \local_node[16].data_out[6] , \local_node[16].data_out[5] , 
        \local_node[16].data_out[4] , \local_node[16].data_out[3] , 
        \local_node[16].data_out[2] , \local_node[16].data_out[1] , 
        \local_node[16].data_out[0] }), .\node_0.clk (\clk.clk ), 
        .\node_0.buffer_full_in (1'b0), .\node_0.receiving_data (1'b0), 
        .\node_0.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_1.clk (
        \clk.clk ), .\node_1.buffer_full_in (1'b0), .\node_1.receiving_data (
        1'b0), .\node_1.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  node4_NODE_X1_NODE_Y0I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__I_node_2_node_interface__ t1 ( 
        .\clk.clk (\clk.clk ), .\reset.reset (\reset.reset ), 
        .\local_node.clk (\local_node[1].clk ), .\local_node.buffer_full_in (
        \local_node[1].buffer_full_in ), .\local_node.buffer_full_out (
        \local_node[1].buffer_full_out ), .\local_node.receiving_data (
        \local_node[1].receiving_data ), .\local_node.sending_data (
        \local_node[1].sending_data ), .\local_node.data_in ({
        \local_node[1].data_in  [15], \local_node[1].data_in  [14], 
        \local_node[1].data_in  [13], \local_node[1].data_in  [12], 
        \local_node[1].data_in  [11], \local_node[1].data_in  [10], 
        \local_node[1].data_in  [9], \local_node[1].data_in  [8], 
        \local_node[1].data_in  [7], \local_node[1].data_in  [6], 
        \local_node[1].data_in  [5], \local_node[1].data_in  [4], 
        \local_node[1].data_in  [3], \local_node[1].data_in  [2], 
        \local_node[1].data_in  [1], \local_node[1].data_in  [0]}), 
        .\local_node.data_out ({\local_node[1].data_out  [15], 
        \local_node[1].data_out  [14], \local_node[1].data_out  [13], 
        \local_node[1].data_out  [12], \local_node[1].data_out  [11], 
        \local_node[1].data_out  [10], \local_node[1].data_out  [9], 
        \local_node[1].data_out  [8], \local_node[1].data_out  [7], 
        \local_node[1].data_out  [6], \local_node[1].data_out  [5], 
        \local_node[1].data_out  [4], \local_node[1].data_out  [3], 
        \local_node[1].data_out  [2], \local_node[1].data_out  [1], 
        \local_node[1].data_out  [0]}), .\node_0.clk (\clk.clk ), 
        .\node_0.buffer_full_in (1'b0), .\node_0.receiving_data (1'b0), 
        .\node_0.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_1.clk (
        \clk.clk ), .\node_1.buffer_full_in (1'b0), .\node_1.receiving_data (
        1'b0), .\node_1.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_2.clk (
        \clk.clk ), .\node_2.buffer_full_in (1'b0), .\node_2.receiving_data (
        1'b0), .\node_2.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  node4_NODE_X2_NODE_Y0I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__I_node_2_node_interface__ t2 ( 
        .\clk.clk (\clk.clk ), .\reset.reset (\reset.reset ), 
        .\local_node.clk (\local_node[2].clk ), .\local_node.buffer_full_in (
        \local_node[2].buffer_full_in ), .\local_node.buffer_full_out (
        \local_node[2].buffer_full_out ), .\local_node.receiving_data (
        \local_node[2].receiving_data ), .\local_node.sending_data (
        \local_node[2].sending_data ), .\local_node.data_in ({
        \local_node[2].data_in  [15], \local_node[2].data_in  [14], 
        \local_node[2].data_in  [13], \local_node[2].data_in  [12], 
        \local_node[2].data_in  [11], \local_node[2].data_in  [10], 
        \local_node[2].data_in  [9], \local_node[2].data_in  [8], 
        \local_node[2].data_in  [7], \local_node[2].data_in  [6], 
        \local_node[2].data_in  [5], \local_node[2].data_in  [4], 
        \local_node[2].data_in  [3], \local_node[2].data_in  [2], 
        \local_node[2].data_in  [1], \local_node[2].data_in  [0]}), 
        .\local_node.data_out ({\local_node[2].data_out  [15], 
        \local_node[2].data_out  [14], \local_node[2].data_out  [13], 
        \local_node[2].data_out  [12], \local_node[2].data_out  [11], 
        \local_node[2].data_out  [10], \local_node[2].data_out  [9], 
        \local_node[2].data_out  [8], \local_node[2].data_out  [7], 
        \local_node[2].data_out  [6], \local_node[2].data_out  [5], 
        \local_node[2].data_out  [4], \local_node[2].data_out  [3], 
        \local_node[2].data_out  [2], \local_node[2].data_out  [1], 
        \local_node[2].data_out  [0]}), .\node_0.clk (\clk.clk ), 
        .\node_0.buffer_full_in (1'b0), .\node_0.receiving_data (1'b0), 
        .\node_0.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_1.clk (
        \clk.clk ), .\node_1.buffer_full_in (1'b0), .\node_1.receiving_data (
        1'b0), .\node_1.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_2.clk (
        \clk.clk ), .\node_2.buffer_full_in (1'b0), .\node_2.receiving_data (
        1'b0), .\node_2.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  node4_NODE_X1_NODE_Y3I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__I_node_2_node_interface__ b1 ( 
        .\clk.clk (\clk.clk ), .\reset.reset (\reset.reset ), 
        .\local_node.clk (\local_node[13].clk ), .\local_node.buffer_full_in (
        \local_node[13].buffer_full_in ), .\local_node.buffer_full_out (
        \local_node[13].buffer_full_out ), .\local_node.receiving_data (
        \local_node[13].receiving_data ), .\local_node.sending_data (
        \local_node[13].sending_data ), .\local_node.data_in ({
        \local_node[13].data_in  [15], \local_node[13].data_in  [14], 
        \local_node[13].data_in  [13], \local_node[13].data_in  [12], 
        \local_node[13].data_in  [11], \local_node[13].data_in  [10], 
        \local_node[13].data_in  [9], \local_node[13].data_in  [8], 
        \local_node[13].data_in  [7], \local_node[13].data_in  [6], 
        \local_node[13].data_in  [5], \local_node[13].data_in  [4], 
        \local_node[13].data_in  [3], \local_node[13].data_in  [2], 
        \local_node[13].data_in  [1], \local_node[13].data_in  [0]}), 
        .\local_node.data_out ({\local_node[13].data_out  [15], 
        \local_node[13].data_out  [14], \local_node[13].data_out  [13], 
        \local_node[13].data_out  [12], \local_node[13].data_out  [11], 
        \local_node[13].data_out  [10], \local_node[13].data_out  [9], 
        \local_node[13].data_out  [8], \local_node[13].data_out  [7], 
        \local_node[13].data_out  [6], \local_node[13].data_out  [5], 
        \local_node[13].data_out  [4], \local_node[13].data_out  [3], 
        \local_node[13].data_out  [2], \local_node[13].data_out  [1], 
        \local_node[13].data_out  [0]}), .\node_0.clk (\clk.clk ), 
        .\node_0.buffer_full_in (1'b0), .\node_0.receiving_data (1'b0), 
        .\node_0.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_1.clk (
        \clk.clk ), .\node_1.buffer_full_in (1'b0), .\node_1.receiving_data (
        1'b0), .\node_1.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_2.clk (
        \clk.clk ), .\node_2.buffer_full_in (1'b0), .\node_2.receiving_data (
        1'b0), .\node_2.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  node4_NODE_X2_NODE_Y3I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__I_node_2_node_interface__ b2 ( 
        .\clk.clk (\clk.clk ), .\reset.reset (\reset.reset ), 
        .\local_node.clk (\local_node[14].clk ), .\local_node.buffer_full_in (
        \local_node[14].buffer_full_in ), .\local_node.buffer_full_out (
        \local_node[14].buffer_full_out ), .\local_node.receiving_data (
        \local_node[14].receiving_data ), .\local_node.sending_data (
        \local_node[14].sending_data ), .\local_node.data_in ({
        \local_node[14].data_in  [15], \local_node[14].data_in  [14], 
        \local_node[14].data_in  [13], \local_node[14].data_in  [12], 
        \local_node[14].data_in  [11], \local_node[14].data_in  [10], 
        \local_node[14].data_in  [9], \local_node[14].data_in  [8], 
        \local_node[14].data_in  [7], \local_node[14].data_in  [6], 
        \local_node[14].data_in  [5], \local_node[14].data_in  [4], 
        \local_node[14].data_in  [3], \local_node[14].data_in  [2], 
        \local_node[14].data_in  [1], \local_node[14].data_in  [0]}), 
        .\local_node.data_out ({\local_node[14].data_out  [15], 
        \local_node[14].data_out  [14], \local_node[14].data_out  [13], 
        \local_node[14].data_out  [12], \local_node[14].data_out  [11], 
        \local_node[14].data_out  [10], \local_node[14].data_out  [9], 
        \local_node[14].data_out  [8], \local_node[14].data_out  [7], 
        \local_node[14].data_out  [6], \local_node[14].data_out  [5], 
        \local_node[14].data_out  [4], \local_node[14].data_out  [3], 
        \local_node[14].data_out  [2], \local_node[14].data_out  [1], 
        \local_node[14].data_out  [0]}), .\node_0.clk (\clk.clk ), 
        .\node_0.buffer_full_in (1'b0), .\node_0.receiving_data (1'b0), 
        .\node_0.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_1.clk (
        \clk.clk ), .\node_1.buffer_full_in (1'b0), .\node_1.receiving_data (
        1'b0), .\node_1.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_2.clk (
        \clk.clk ), .\node_2.buffer_full_in (1'b0), .\node_2.receiving_data (
        1'b0), .\node_2.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  node4_NODE_X0_NODE_Y1I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__I_node_2_node_interface__ l1 ( 
        .\clk.clk (\clk.clk ), .\reset.reset (\reset.reset ), 
        .\local_node.clk (\local_node[4].clk ), .\local_node.buffer_full_in (
        \local_node[4].buffer_full_in ), .\local_node.buffer_full_out (
        \local_node[4].buffer_full_out ), .\local_node.receiving_data (
        \local_node[4].receiving_data ), .\local_node.sending_data (
        \local_node[4].sending_data ), .\local_node.data_in ({
        \local_node[4].data_in  [15], \local_node[4].data_in  [14], 
        \local_node[4].data_in  [13], \local_node[4].data_in  [12], 
        \local_node[4].data_in  [11], \local_node[4].data_in  [10], 
        \local_node[4].data_in  [9], \local_node[4].data_in  [8], 
        \local_node[4].data_in  [7], \local_node[4].data_in  [6], 
        \local_node[4].data_in  [5], \local_node[4].data_in  [4], 
        \local_node[4].data_in  [3], \local_node[4].data_in  [2], 
        \local_node[4].data_in  [1], \local_node[4].data_in  [0]}), 
        .\local_node.data_out ({\local_node[4].data_out  [15], 
        \local_node[4].data_out  [14], \local_node[4].data_out  [13], 
        \local_node[4].data_out  [12], \local_node[4].data_out  [11], 
        \local_node[4].data_out  [10], \local_node[4].data_out  [9], 
        \local_node[4].data_out  [8], \local_node[4].data_out  [7], 
        \local_node[4].data_out  [6], \local_node[4].data_out  [5], 
        \local_node[4].data_out  [4], \local_node[4].data_out  [3], 
        \local_node[4].data_out  [2], \local_node[4].data_out  [1], 
        \local_node[4].data_out  [0]}), .\node_0.clk (\clk.clk ), 
        .\node_0.buffer_full_in (1'b0), .\node_0.receiving_data (1'b0), 
        .\node_0.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_1.clk (
        \clk.clk ), .\node_1.buffer_full_in (1'b0), .\node_1.receiving_data (
        1'b0), .\node_1.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_2.clk (
        \clk.clk ), .\node_2.buffer_full_in (1'b0), .\node_2.receiving_data (
        1'b0), .\node_2.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  node4_NODE_X0_NODE_Y2I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__I_node_2_node_interface__ l2 ( 
        .\clk.clk (\clk.clk ), .\reset.reset (\reset.reset ), 
        .\local_node.clk (\local_node[8].clk ), .\local_node.buffer_full_in (
        \local_node[8].buffer_full_in ), .\local_node.buffer_full_out (
        \local_node[8].buffer_full_out ), .\local_node.receiving_data (
        \local_node[8].receiving_data ), .\local_node.sending_data (
        \local_node[8].sending_data ), .\local_node.data_in ({
        \local_node[8].data_in  [15], \local_node[8].data_in  [14], 
        \local_node[8].data_in  [13], \local_node[8].data_in  [12], 
        \local_node[8].data_in  [11], \local_node[8].data_in  [10], 
        \local_node[8].data_in  [9], \local_node[8].data_in  [8], 
        \local_node[8].data_in  [7], \local_node[8].data_in  [6], 
        \local_node[8].data_in  [5], \local_node[8].data_in  [4], 
        \local_node[8].data_in  [3], \local_node[8].data_in  [2], 
        \local_node[8].data_in  [1], \local_node[8].data_in  [0]}), 
        .\local_node.data_out ({\local_node[8].data_out  [15], 
        \local_node[8].data_out  [14], \local_node[8].data_out  [13], 
        \local_node[8].data_out  [12], \local_node[8].data_out  [11], 
        \local_node[8].data_out  [10], \local_node[8].data_out  [9], 
        \local_node[8].data_out  [8], \local_node[8].data_out  [7], 
        \local_node[8].data_out  [6], \local_node[8].data_out  [5], 
        \local_node[8].data_out  [4], \local_node[8].data_out  [3], 
        \local_node[8].data_out  [2], \local_node[8].data_out  [1], 
        \local_node[8].data_out  [0]}), .\node_0.clk (\clk.clk ), 
        .\node_0.buffer_full_in (1'b0), .\node_0.receiving_data (1'b0), 
        .\node_0.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_1.clk (
        \clk.clk ), .\node_1.buffer_full_in (1'b0), .\node_1.receiving_data (
        1'b0), .\node_1.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_2.clk (
        \clk.clk ), .\node_2.buffer_full_in (1'b0), .\node_2.receiving_data (
        1'b0), .\node_2.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  node4_NODE_X3_NODE_Y1I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__I_node_2_node_interface__ r1 ( 
        .\clk.clk (\clk.clk ), .\reset.reset (\reset.reset ), 
        .\local_node.clk (\local_node[7].clk ), .\local_node.buffer_full_in (
        \local_node[7].buffer_full_in ), .\local_node.buffer_full_out (
        \local_node[7].buffer_full_out ), .\local_node.receiving_data (
        \local_node[7].receiving_data ), .\local_node.sending_data (
        \local_node[7].sending_data ), .\local_node.data_in ({
        \local_node[7].data_in  [15], \local_node[7].data_in  [14], 
        \local_node[7].data_in  [13], \local_node[7].data_in  [12], 
        \local_node[7].data_in  [11], \local_node[7].data_in  [10], 
        \local_node[7].data_in  [9], \local_node[7].data_in  [8], 
        \local_node[7].data_in  [7], \local_node[7].data_in  [6], 
        \local_node[7].data_in  [5], \local_node[7].data_in  [4], 
        \local_node[7].data_in  [3], \local_node[7].data_in  [2], 
        \local_node[7].data_in  [1], \local_node[7].data_in  [0]}), 
        .\local_node.data_out ({\local_node[7].data_out  [15], 
        \local_node[7].data_out  [14], \local_node[7].data_out  [13], 
        \local_node[7].data_out  [12], \local_node[7].data_out  [11], 
        \local_node[7].data_out  [10], \local_node[7].data_out  [9], 
        \local_node[7].data_out  [8], \local_node[7].data_out  [7], 
        \local_node[7].data_out  [6], \local_node[7].data_out  [5], 
        \local_node[7].data_out  [4], \local_node[7].data_out  [3], 
        \local_node[7].data_out  [2], \local_node[7].data_out  [1], 
        \local_node[7].data_out  [0]}), .\node_0.clk (\clk.clk ), 
        .\node_0.buffer_full_in (1'b0), .\node_0.receiving_data (1'b0), 
        .\node_0.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_1.clk (
        \clk.clk ), .\node_1.buffer_full_in (1'b0), .\node_1.receiving_data (
        1'b0), .\node_1.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_2.clk (
        \clk.clk ), .\node_2.buffer_full_in (1'b0), .\node_2.receiving_data (
        1'b0), .\node_2.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  node4_NODE_X3_NODE_Y2I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__I_node_2_node_interface__ r2 ( 
        .\clk.clk (\clk.clk ), .\reset.reset (\reset.reset ), 
        .\local_node.clk (\local_node[11].clk ), .\local_node.buffer_full_in (
        \local_node[11].buffer_full_in ), .\local_node.buffer_full_out (
        \local_node[11].buffer_full_out ), .\local_node.receiving_data (
        \local_node[11].receiving_data ), .\local_node.sending_data (
        \local_node[11].sending_data ), .\local_node.data_in ({
        \local_node[11].data_in  [15], \local_node[11].data_in  [14], 
        \local_node[11].data_in  [13], \local_node[11].data_in  [12], 
        \local_node[11].data_in  [11], \local_node[11].data_in  [10], 
        \local_node[11].data_in  [9], \local_node[11].data_in  [8], 
        \local_node[11].data_in  [7], \local_node[11].data_in  [6], 
        \local_node[11].data_in  [5], \local_node[11].data_in  [4], 
        \local_node[11].data_in  [3], \local_node[11].data_in  [2], 
        \local_node[11].data_in  [1], \local_node[11].data_in  [0]}), 
        .\local_node.data_out ({\local_node[11].data_out  [15], 
        \local_node[11].data_out  [14], \local_node[11].data_out  [13], 
        \local_node[11].data_out  [12], \local_node[11].data_out  [11], 
        \local_node[11].data_out  [10], \local_node[11].data_out  [9], 
        \local_node[11].data_out  [8], \local_node[11].data_out  [7], 
        \local_node[11].data_out  [6], \local_node[11].data_out  [5], 
        \local_node[11].data_out  [4], \local_node[11].data_out  [3], 
        \local_node[11].data_out  [2], \local_node[11].data_out  [1], 
        \local_node[11].data_out  [0]}), .\node_0.clk (\clk.clk ), 
        .\node_0.buffer_full_in (1'b0), .\node_0.receiving_data (1'b0), 
        .\node_0.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_1.clk (
        \clk.clk ), .\node_1.buffer_full_in (1'b0), .\node_1.receiving_data (
        1'b0), .\node_1.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_2.clk (
        \clk.clk ), .\node_2.buffer_full_in (1'b0), .\node_2.receiving_data (
        1'b0), .\node_2.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  node5_NODE_X1_NODE_Y1I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__I_node_2_node_interface__I_node_3_node_interface__ n1 ( 
        .\clk.clk (\clk.clk ), .\reset.reset (\reset.reset ), 
        .\local_node.clk (\local_node[5].clk ), .\local_node.buffer_full_in (
        \local_node[5].buffer_full_in ), .\local_node.buffer_full_out (
        \local_node[5].buffer_full_out ), .\local_node.receiving_data (
        \local_node[5].receiving_data ), .\local_node.sending_data (
        \local_node[5].sending_data ), .\local_node.data_in ({
        \local_node[5].data_in  [15], \local_node[5].data_in  [14], 
        \local_node[5].data_in  [13], \local_node[5].data_in  [12], 
        \local_node[5].data_in  [11], \local_node[5].data_in  [10], 
        \local_node[5].data_in  [9], \local_node[5].data_in  [8], 
        \local_node[5].data_in  [7], \local_node[5].data_in  [6], 
        \local_node[5].data_in  [5], \local_node[5].data_in  [4], 
        \local_node[5].data_in  [3], \local_node[5].data_in  [2], 
        \local_node[5].data_in  [1], \local_node[5].data_in  [0]}), 
        .\local_node.data_out ({\local_node[5].data_out  [15], 
        \local_node[5].data_out  [14], \local_node[5].data_out  [13], 
        \local_node[5].data_out  [12], \local_node[5].data_out  [11], 
        \local_node[5].data_out  [10], \local_node[5].data_out  [9], 
        \local_node[5].data_out  [8], \local_node[5].data_out  [7], 
        \local_node[5].data_out  [6], \local_node[5].data_out  [5], 
        \local_node[5].data_out  [4], \local_node[5].data_out  [3], 
        \local_node[5].data_out  [2], \local_node[5].data_out  [1], 
        \local_node[5].data_out  [0]}), .\node_0.clk (\clk.clk ), 
        .\node_0.buffer_full_in (1'b0), .\node_0.receiving_data (1'b0), 
        .\node_0.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_1.clk (
        \clk.clk ), .\node_1.buffer_full_in (1'b0), .\node_1.receiving_data (
        1'b0), .\node_1.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_2.clk (
        \clk.clk ), .\node_2.buffer_full_in (1'b0), .\node_2.receiving_data (
        1'b0), .\node_2.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_3.clk (
        \clk.clk ), .\node_3.buffer_full_in (1'b0), .\node_3.receiving_data (
        1'b0), .\node_3.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  node5_NODE_X1_NODE_Y2I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__I_node_2_node_interface__I_node_3_node_interface__ n2 ( 
        .\clk.clk (\clk.clk ), .\reset.reset (\reset.reset ), 
        .\local_node.clk (\local_node[9].clk ), .\local_node.buffer_full_in (
        \local_node[9].buffer_full_in ), .\local_node.buffer_full_out (
        \local_node[9].buffer_full_out ), .\local_node.receiving_data (
        \local_node[9].receiving_data ), .\local_node.sending_data (
        \local_node[9].sending_data ), .\local_node.data_in ({
        \local_node[9].data_in  [15], \local_node[9].data_in  [14], 
        \local_node[9].data_in  [13], \local_node[9].data_in  [12], 
        \local_node[9].data_in  [11], \local_node[9].data_in  [10], 
        \local_node[9].data_in  [9], \local_node[9].data_in  [8], 
        \local_node[9].data_in  [7], \local_node[9].data_in  [6], 
        \local_node[9].data_in  [5], \local_node[9].data_in  [4], 
        \local_node[9].data_in  [3], \local_node[9].data_in  [2], 
        \local_node[9].data_in  [1], \local_node[9].data_in  [0]}), 
        .\local_node.data_out ({\local_node[9].data_out  [15], 
        \local_node[9].data_out  [14], \local_node[9].data_out  [13], 
        \local_node[9].data_out  [12], \local_node[9].data_out  [11], 
        \local_node[9].data_out  [10], \local_node[9].data_out  [9], 
        \local_node[9].data_out  [8], \local_node[9].data_out  [7], 
        \local_node[9].data_out  [6], \local_node[9].data_out  [5], 
        \local_node[9].data_out  [4], \local_node[9].data_out  [3], 
        \local_node[9].data_out  [2], \local_node[9].data_out  [1], 
        \local_node[9].data_out  [0]}), .\node_0.clk (\clk.clk ), 
        .\node_0.buffer_full_in (1'b0), .\node_0.receiving_data (1'b0), 
        .\node_0.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_1.clk (
        \clk.clk ), .\node_1.buffer_full_in (1'b0), .\node_1.receiving_data (
        1'b0), .\node_1.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_2.clk (
        \clk.clk ), .\node_2.buffer_full_in (1'b0), .\node_2.receiving_data (
        1'b0), .\node_2.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_3.clk (
        \clk.clk ), .\node_3.buffer_full_in (1'b0), .\node_3.receiving_data (
        1'b0), .\node_3.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  node5_NODE_X2_NODE_Y1I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__I_node_2_node_interface__I_node_3_node_interface__ n3 ( 
        .\clk.clk (\clk.clk ), .\reset.reset (\reset.reset ), 
        .\local_node.clk (\local_node[6].clk ), .\local_node.buffer_full_in (
        \local_node[6].buffer_full_in ), .\local_node.buffer_full_out (
        \local_node[6].buffer_full_out ), .\local_node.receiving_data (
        \local_node[6].receiving_data ), .\local_node.sending_data (
        \local_node[6].sending_data ), .\local_node.data_in ({
        \local_node[6].data_in  [15], \local_node[6].data_in  [14], 
        \local_node[6].data_in  [13], \local_node[6].data_in  [12], 
        \local_node[6].data_in  [11], \local_node[6].data_in  [10], 
        \local_node[6].data_in  [9], \local_node[6].data_in  [8], 
        \local_node[6].data_in  [7], \local_node[6].data_in  [6], 
        \local_node[6].data_in  [5], \local_node[6].data_in  [4], 
        \local_node[6].data_in  [3], \local_node[6].data_in  [2], 
        \local_node[6].data_in  [1], \local_node[6].data_in  [0]}), 
        .\local_node.data_out ({\local_node[6].data_out  [15], 
        \local_node[6].data_out  [14], \local_node[6].data_out  [13], 
        \local_node[6].data_out  [12], \local_node[6].data_out  [11], 
        \local_node[6].data_out  [10], \local_node[6].data_out  [9], 
        \local_node[6].data_out  [8], \local_node[6].data_out  [7], 
        \local_node[6].data_out  [6], \local_node[6].data_out  [5], 
        \local_node[6].data_out  [4], \local_node[6].data_out  [3], 
        \local_node[6].data_out  [2], \local_node[6].data_out  [1], 
        \local_node[6].data_out  [0]}), .\node_0.clk (\clk.clk ), 
        .\node_0.buffer_full_in (1'b0), .\node_0.receiving_data (1'b0), 
        .\node_0.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_1.clk (
        \clk.clk ), .\node_1.buffer_full_in (1'b0), .\node_1.receiving_data (
        1'b0), .\node_1.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_2.clk (
        \clk.clk ), .\node_2.buffer_full_in (1'b0), .\node_2.receiving_data (
        1'b0), .\node_2.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_3.clk (
        \clk.clk ), .\node_3.buffer_full_in (1'b0), .\node_3.receiving_data (
        1'b0), .\node_3.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  node5_NODE_X2_NODE_Y2I_clk_clock_interface_dut_I_reset_reset_interface_dut_I_local_node_node_interface__I_node_0_node_interface__I_node_1_node_interface__I_node_2_node_interface__I_node_3_node_interface__ n4 ( 
        .\clk.clk (\clk.clk ), .\reset.reset (\reset.reset ), 
        .\local_node.clk (\local_node[10].clk ), .\local_node.buffer_full_in (
        \local_node[10].buffer_full_in ), .\local_node.buffer_full_out (
        \local_node[10].buffer_full_out ), .\local_node.receiving_data (
        \local_node[10].receiving_data ), .\local_node.sending_data (
        \local_node[10].sending_data ), .\local_node.data_in ({
        \local_node[10].data_in  [15], \local_node[10].data_in  [14], 
        \local_node[10].data_in  [13], \local_node[10].data_in  [12], 
        \local_node[10].data_in  [11], \local_node[10].data_in  [10], 
        \local_node[10].data_in  [9], \local_node[10].data_in  [8], 
        \local_node[10].data_in  [7], \local_node[10].data_in  [6], 
        \local_node[10].data_in  [5], \local_node[10].data_in  [4], 
        \local_node[10].data_in  [3], \local_node[10].data_in  [2], 
        \local_node[10].data_in  [1], \local_node[10].data_in  [0]}), 
        .\local_node.data_out ({\local_node[10].data_out  [15], 
        \local_node[10].data_out  [14], \local_node[10].data_out  [13], 
        \local_node[10].data_out  [12], \local_node[10].data_out  [11], 
        \local_node[10].data_out  [10], \local_node[10].data_out  [9], 
        \local_node[10].data_out  [8], \local_node[10].data_out  [7], 
        \local_node[10].data_out  [6], \local_node[10].data_out  [5], 
        \local_node[10].data_out  [4], \local_node[10].data_out  [3], 
        \local_node[10].data_out  [2], \local_node[10].data_out  [1], 
        \local_node[10].data_out  [0]}), .\node_0.clk (\clk.clk ), 
        .\node_0.buffer_full_in (1'b0), .\node_0.receiving_data (1'b0), 
        .\node_0.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_1.clk (
        \clk.clk ), .\node_1.buffer_full_in (1'b0), .\node_1.receiving_data (
        1'b0), .\node_1.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_2.clk (
        \clk.clk ), .\node_2.buffer_full_in (1'b0), .\node_2.receiving_data (
        1'b0), .\node_2.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\node_3.clk (
        \clk.clk ), .\node_3.buffer_full_in (1'b0), .\node_3.receiving_data (
        1'b0), .\node_3.data_in ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
endmodule

