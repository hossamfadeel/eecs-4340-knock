class data;
endclass
