module node4(
	clk_interface.dut clk,
	reset_interface.dut reset,
	node_interface.dut local_node,
	node_interface.dut node_0,
	node_interface.dut node_1,
	node_interface.dut node_2
);


endmodule
