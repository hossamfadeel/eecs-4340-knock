`define TOP(y) y==0
`define BOTTOM(y) y==`NOC_SIZE
`define LEFT(x) x==0
`define RIGHT(x) x==`NOC_SIZE
