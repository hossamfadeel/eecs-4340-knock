`define NSMO (`NOC_SIZE-1) 

`define TOP(y) y==0
`define BOTTOM(y) y==`NSMO
`define LEFT(x) x==0
`define RIGHT(x) x==`NSMO
