class environment;
  data d;
  configuration cfg;
  tracker t;
  reset_transaction rst;

  function new();
    d = new();
    cfg = new();
    t = new();

    rst = new(this);
  endfunction

  function gen();

  endfunction

  function check();

  endfunction

  function shift();

  endfunction
endclass
